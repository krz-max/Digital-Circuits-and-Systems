//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ChvCTq9WgOpXAwrNAcHqo3WDy8IEdM/HHpU8e2J+TqSnizttBYxqyKJpDoROKAMv
CQ76E+3GUCI4UaCvl7YjSZDVgXJNCD743sdqboYcrULc0iB6h+qqKjZ1MYRvmK+l
XJriXcMR769EF2C3YXJt9zgqMzBKmAd8tTEwmOyYL3jx/Q2J3v4Isg==
//pragma protect end_key_block
//pragma protect digest_block
rcdhNwWkc6CmdWGW3T1Ttab6b9U=
//pragma protect end_digest_block
//pragma protect data_block
Dwe4dD9v0h63FkvF4/H8yga/TR01mwTdo+XJQRqIeW9Closm5pqGeVOfW3FAxpIt
a4B3xKAyoFvMrGxZQ+RQQtKaa/qlcslSQDEJZ/tTCKQXAcyUPorLXk9xiLEe2xuR
bIx3hCRNiTN1Ni4C5NHhGWJqfpYN0xYsb29dvrt9KR9sqL4wlmuYkJx+O/oxfkp8
20aab92uriEpROGpaRKIZxHRV1qZsbGQrAC1fOI4KwW7wvx+ZWXxU/4Az7dgXkuf
xUIOH1Xx4Zu6/GqNiCPIlCZSYYBHGv1z1W72LcEJu+SottFtYk46u0zuPqCFmmJD
ow1KrHODnU9IQJ5bRhpD6kVmU32qLm8aEkyKeXabEsVN5F0jfD/ry6eQxxjjpWtI
XECL7zB/hej53PVPBmIHMsPyl1FAYGr4fdrGYDOCdrngYiS5v+YWT8Io5YIjtL7S
uzTrFu06kv3RqKi8nB37dJn4n+QbFJbfxEQd29jx/a/U0/IwvapUnUfYRZswpbM5
b6IuouVCF5g9Bef9Ie5WaOzmX5TcoCU/zdGDSPPdSMvHdRHN+dJdl9EMHJL0OTuD
eldcflOp4fK3DTcUPp2Iy8dFN1lqPsonNb6xZAJsAQr1CyrUbf6BbJKKrkAXu6Ds
dDv9KFm2hJehwh8aqrjH9ksL/EvDeqeScV5QBArt4sPB61LPTJEiudRDfYTHW1fx
mr+uqFxGv7CRVg5Iee9DTjGhgZu33oXbkS8Rs0IlMYw11JmlFAVWKy2munwrRkyZ
c9aL3CkKvZ4aYOdWjIr6f3jKtSyDMNW+Zwp5hJVR2yv5QcyPkgb6nfXp3tH1JlKi
Z33a0dqRa2WCdca0tcidxc4UcvUPPG6mtcTpVQzv/6I0r8OZP8woyl5/e7TFCPdr
HtP3QsHN1sDH9EP6s4sUeaaBgGaiHtl4uCRcnAHcPzpvNd5uGHxvAmhiBRJG9N9P
5oyhWhvf+jt3UVI+yh86bfYqZFs0Nv1zCRLHJ+HW89qn8SbZSWvRQ5fvSKT56plX
MijxI5DypuFhbGjIJtVqrT7/Ba7KaOKh5cIsRO+AIgcLhAx+vzgjD/VCrI7aagUV
Wfx9q+8UYn1tC59CeVDJz3Rp1c4JemsgeqahQ3DTcXsXqWRsgbsvBTZnATGJ6i3M
609cMeETn8n1TyC0tywULTsXi1GV7/AzjCnqEFCkFV5bhrcpdsaQztarDMn+nsH+
Y7WCr34LLWc0KKuoHx+Z66ATMfzDscpsaWTM9Ec7+Ow3bzwQW5WP59YSNOhg8s+P
k2FYqeFWtJLSdku4wPgtGdU9IKxe1+KgMUSIh0OKrSOzd/+jQHNqj6CddrvXJFmi
mU82vGS2ZB7/7KhbHGKt2RsVR59SJG7eF2pXuuT8OEiyrvDZNLfyLvyPgoGYooUJ
LGpptPJ4d7J6Spc3VlglhjZ6tXG3b7VNJmaPfXk1vzA8B7AulgyzDaX0v/OcTraI
Be+nSyE+r1FmtjH362RtYQRcc/Z1Y1RaxWKeeSLR20jIyNSLznxGMaaCOITAobdh
ox8e3X8iA9namajS9n1bkZkk2uGYB3QWrJPRnWNdlDh1LD0OGIgogNKFddeDsNa8
xQdfERoxoFww3WC+FQrxirlKoY/zLECWBSYrYPI2Qu5VnMMhN9Dnzaqn7sg7PgNI
hrb9S88Q6yTvMnAAxUIK2RPWMFzMbT2AqWGlsz0Z/h4OYOds2+pqpUX0cusVZnr6
KJjSQxxvY/Up0EDhQ7fiYLvselhq2+z3jzek/pVJo5oIX5CeBN32odb5gcG/DfoA
X7rk9XJqM5j6IrSG5ePbpciRec0qDjo5El/I9GYWROnzDDSfElbTA1ng+bC7MYqD
MMygy9q9AMT+hdeV7f4G6p6OIR1vMj5Z2bMRbWC6YNK7DHViR/odr4Q70QUFlvk0
aEeL3K5T6/UofqMDLBYQwttsMArPMGz5RQpwfDFQdfj7OajsZnjQCSksiOkNxtNj
XSer9IwPEmGHKQdkb9wienr1IHAQ9Zh+GQfhxrFpHQhLcQSBFe2Q5rYWmxG9qIBG
RIoaHDX68xhCQJyexcYkboreneNkH3yJsYXjdxiuNVpVX6J572Ffxy1LfiRS8+Tv
9LR4tXbX8zwtQOpZ9nidCgE+cSccBkOelJhkjpeQ6EPy98JE2pM8jREL4RcR31aL
Vtg0SZN6H0gSK0DCTgUKfrlblj+2LV7XnAAGYY4JilNsYoH5popMeZAs9cvz5yYe
WjFs3nYL1sDgLOQ59g/DOCKcHAaTs6RBzmNDzXWgizYLgud4Np8tg0o+iWShOi01
qUi3kJyEmOoJ9wWU0KqTDwqOLy8nL+uXETtNwgmH5U7aKWBgBhg1ME5b+0b+EaDF
R/g74j1wov+gIGUHqqXy5BhzFQEYjPVrGkkJnSS105a7zbqZR53Lctv/6xMzjlGn
9H6GpDWozTTuDfwFjFTtehgI3JizDIMi6E9X8VLxh/uIdKZKyaegYhchAis8rh95
TKiU3jdSdjpWExFSu22YTVxj6nBtpd2dnKnGIkbJEvj5bNU+kg1b94Lm8eWBW6XX
Q1dICpEsYZG7OZDwIgaFWWw0AcJXch2qheopKE7E0Fibs+06SxB6EgfLq1cXh8jb
CZT/777V2H4Zhcywj2H8NRToNpaZwXKu5rwrh7OKaPTCH0YDLj+40Wol7X/2KLGT
JcPYmgEFH61E5E8gJA+2IqzN5ZE2Ilo4r8saxEcl5OXCc+IOYJtFaaMaQkcF77t4
icUO1eDRj9/oDqYSzgVg1qlhhEB5p9br2OjKt3DoZmj2htNYeojGHQYZXcFNgaX3
wAT/zijw1Sq8xSkGgBJgrHL9rkVxRudpkGOGxxj1dLpioHUBHe5B5LxQ7MVAoyxg
1wsZ4i5yaBCNfpRavigqQ7Ns/QY62QHknO/+M6nHlpAZHoS6gBuhSwFZSPNVTKFh
Et3u273/S8opHUzdrKoVQoVVfb+NbPD7JpS4+wt0wh6dHyRCTa5jH560WEhmgcvi
DaIUEUq+icTLpbIj6mTWV8K2Wka+Sxx507ZMZHb3LYHaltsvH6UalxGA3TOUm3tf
FFoGdFLYB0TWSR7ISX+5AGPRMetVTJakv+1v0bGz7VdFX4XvQ096T8KkRkIWCXr/
k7nZLLLwize5MSF2TL6ETvqqhwSUs+hE7O0nKR/ETIncYxp0AoLkaV4AJMIjOv4c
XkeelXyioTFCA9MoJQq7fQiHENTFpcoPTEu2Jfkjox7QN6OMvlYD+959dOy1DRml
iUQB6lruo/51tsKsRkT9F+q86soXFQa6ayKAx+zB6eUZkRGGvr3OvnSPEwfgtVKl
gELx1Cf+BZg7QTZVDhjcjNPpbJd+2VkHrav0wZCkWMV0RIsZrXja0vHWfP+renci
8bVGGZqbUbRTSqE53Q+a9aUipNhAIqFpdsWuQr1cP+7D4ZW3elOKBlz0FOykJbVy
/gf1F/md4tOrPEVnkVoq0H0z5rbOullxNbEy/lkoBo1XHBXDBdU60XQ1cD6OJVgj
o7iOwHA/hB8yxw9EcW3XLVa798lWtuTGvc8dS4CjbdK7ZAaQHr03hml0VPLPK4DW
0Agc0c8QRGU+rln9NUDwi84PdGqPDkhGtfwm2ilwQKptJz4r3FggEaUE9zdwIVG2
xZO1O9cymdqaWCARNOfmB/gQvhtcpc5beNEjcPmfXPzSg/DTdrBldM13ZWwktqXI
ipwp1fbl0/5ngkPzhk+fi6D8YWBRsxblIqbXa4tvuheBXCixpWjS1U6GLzpXPBkw
4zq0alVN+3kPazDRyTDjhVx5xDVs5WHnis5AekqFCqHZVvF8ZUeklHnlkrwcwQ0M
+jJuCoo9gsVGJLTAx/GccgoEC9BkKTJfV0JooQrtLIYZgW2rdOcJnpfTda9a0lKr
09Bw/TCrQwmBgaFK2NmLI1+I7w0GUeL/VqACjuZ9Ypg8i7/W0AO/SNt7S8fSCgO0
UKm1i+kr6Lp207C3EIwcxMPggIVuYCwj4ymSxbAb2zsRq7iKMYCUp+x0LHib0HKb
lHiw/Yva5gXkAJrZfGWQ0v7HVG6Z+9wWidy6UjCxKaZkvL2IT168tjfFOSxZjvFT
qvBoio5SYShxe/BGWx5Z1L+dA47ql1VY5f0VPvRwShIFvuPN76dXndrGDByTMwy5
3nWh2u/GaWyzhvvD8ZrLEgg1hlaLDNekUjVoUbrNRLUS5Bl++IDXlpnDyCi1JN41
RfwAVxr9tL2Rw1jFqmrHj6Wo8RasiNyEI+PN9Yg3pqwTkGkfpofdgxSzWw6uAWT0
YOv/wl7hzhpv2JpRkm1ydb1ntBgk160uHR/s+0psFNzxWBsIBGwra4hum/M048G4
pZe4wpLmYzEIyuTkuvcpw3+/S8+GinzFoycXU2f4IZEOiANcQYnDyLv6a8lV35ZN
dSXVbY6rC5yWuvY7OhtMpH5Xx1+7gZ3OCcM8EODXfeKykNN9ZU5gkAlF72pPGqaL
nS52G4ygvDFrTI/sbCUQBiJP/cUYH/CopxKpCJT6in4pnP1FkI3rq+rdKV2eqIlH
p3hCT640ex71tBor3hc/Bq0+D9ptHSxJoXY8YmjKH4PB7YrZntcxDxarUWArIrYe
6U/mVVnYHt+h3ouNPHchBFbkvxqbp398jeErqeAdidydsa1PBXylurCbty6rdD3f
kjoqN4OAREc2kSpvzxQg+mu3LYAV/77gB+lYzwGJGV64nfSPq3Wpqv8GKRjVgIkJ
U5cmGhh7BsH9CpJlbxuiaxYcMoDK9jx6Wjn33gqBLhnbZTL3Yl/nv8ihrxb88WvD
JCUZIlWkjOXsSNl7wIiD5t+w8vsZtIY7fujB4KlQxjeK918Xg1wl1GSinUWGFixG
jHz8F4oHVOG5j+o85nwMnIG7pDa1lRaAVKSUuIef2NVYLzi7+f8d7RXY+oTXsSo2
E3HPmkW7XJ7bOqxxBjfNFkjU13QLsbqgt+T9lopkv5MraUhGGaaHEF/9LMNFiJBt
hiDBTOV5+XEqvTWVedh1T84wK1mxSehHTfYQJQDb7QRf7ufdNEVHW5eoeVW1v8V/
CUpPShE454WDBkUV2lrS2y9NbTRNVbotITuGx/CfDjRqcxCF6EqVngpU6YOQQMXN
97L+Zi789QQCgNGdW6RMm2WgAReGQPc0WzopD2+IP+ptmT1qQC4aK6/xMTSFxYCV
4co5yxE2QPnQaxCqXTPTCBSiwYt7yZooohjyfANLyUmxCYnzThc3nFY3b8C5yLOe
PrPruSk+e9k+TarRlsXqEda7K6Onv302lKz2UqezRg9aqnsECsJDRBtQfhzdFHRs
PDKrFmi13xLaby5CnL7qMznOu7vzR2M/ImjGHkBU47fnYSvlK9XlkBkP0DmWXnwX
zPy/olRHbMhQ6DbP6TATfCqRit0nK5VbppusM+MjbeyE0lNjqS40TCJdx5dUn55a
SlZaVD6FcN8gk8r9V4rM3jObmSamVOtP11Qm2MDPu3GZPGYUSZMGlpzhosYx4evR
/etGcAS1FLZoS6tbkKLG/lexZWob2xJtAMo2yVOvsz5scdzaIa0pJpeSo6PH4h3w
G3YEYGlHEJMtdB2tUN5KMV/xBEVAvZy7mfSjSrdAMN34EIjzadAgkPh3S5tk+W6W
KF+7EsNWJUOW+wlSfQT6vuwmbGMsdYGk2/dgvQ6AzIXBEr09LGSBB/EMEz88hUtL
dSwnuI7fMBxi7Lh5lbGND9mcOy4pHnXwbsJ0Zy049jKJU/rZxYtFbDPwjUStm7O5
x8ZLiiN30xHSJ2DbXd7ddXZ2UkJ8GxJsyA6qHFDwXXKnpU9/74S1mjGtoiSy2B/N
GiHnP32Df0xrO1kYf+YyXxCY1I716I5wlz6x1ZN1pXVwioQ+BI90+HpnsWHrXSW2
drAn3zQ7Z2X14xjELEeupAGkTrVvK83H1R93NLsS4DNSiNBHOm4bHbrgD8sfWNYV
vx2eC1F5Mv/qpoI4HbrPdS4AskP4sR5Y4TXF8NcVPA6RzNUuiZeoxe98szQ4azOC
sshHAJYWnJr/qnUqnQfVgfKcp4DQszS7M40/o+qR9GTWGgYbhbnteUHdXnKyGSK6
JyynGD49zJtsWpfJC+SnTaHw4mgYi+rN+GI2MFjR7AhunHuGGmgFitZ2LmiY+OHi
550quR6GZXCA9YTdCmSaYGQsUL2jQuud7W3jTU7h+MU+eCkfJ5cc18C902JFtSkS
ThEMemWzkXRAYtnYraO2I0/dqaeObNQcex+78TeJU0BZ4lPrI5VPiiSt+WA+6ptn
eLnvxMXQkwPbY326X2TDXjY011SCg1s/pke/ZrBtPB6yKykD12vvD8iog8ijnpnp
pwmyYtllpMeOmhO9wiVbrTL1UlzmkLvhbQNZJHPbWKDKwS0LOAtEBgPVCHvAq1JF
7Yl3IY3O9rcniP+W3xV4879cdJAiPNJsdgDLsSW02tP0gwhjYocxFaQqjF4+0TSJ
vr66R0l937k4vi34J1FHKftzu1Vq5v45XT35OF1+GxWJUZvCd+94El97+/QwB5EB
AmOukGU7TEctLerNhQCuYI0/SIAa4WEgFveG10wE0hA02u7+9nZvHx2ZAhLyjuqo
mouBibQxFbq1XAIwPdtI5xN4l0tAWELHgwCidskqTCsgKtw2IIY+0DYBaF4+3njp
JtGxWolj8dznrsVcL2IZCmhi4bVzDiFBWvdGOiivCrmucNGOEev2CA34dIX1smQw
NVysbnT4N/2/4LKv7fruOOQc3iwWCdK9NlCtPNGp21KMP1tp6GmDHZEzZztjvZbk
YjPGyu0LyA9YtEfAXBK+VNEVW4RbgD6PDBEmqUhmRziPYgUK/wH36rV30Dl3SZHH
8OjyF94MNJ+4ioirf/6MaekLpc07WiErtj8CTIeS0R+kKYMMCeIQvMFI8ndwWt7V
0tsNEiMh3GYLwzxm/xsVT8b+2xg2ZYh+OLM959TPyeh972SvE7EvMTWip9Q2g3TU
aMlsLr8QszsEQpziF+JH+/lGFsY76t/wZ/evB8TZf9CgC6Wnsy4FeuoYh7216ujo
XlVujCVWcldMtRkPMxRRCW1PgMUW07ej/xp9XgzU6DVuKLgFtiaWy/KQJL7DofRd
fH/zIrosWc3S/bLas4qPYBAAxRuVadO3+FyC1+9kH5hnU0snG7uU6xxuwp2j2pEx
rVte9WgcmdCwm8zgNoYSUjT7SxJUoOMEByQKqZqIPjBvsdyTPZXUBymgSD8e/YuI
10bMm1JAjZb1n0545hBZbKxo+XsGbVw5u0GXmZxX4ig=
//pragma protect end_data_block
//pragma protect digest_block
rrfkp4hRMciZzhnFQr5E/ju40B0=
//pragma protect end_digest_block
//pragma protect end_protected
