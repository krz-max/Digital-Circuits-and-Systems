//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
oUSHxiTbF4AL7Rt4FeqeWlp/1m/fusDelHEaXxdea2LXLHhD3LQoezxMS84vYHM3
WlZcmYEGHgWCjXXiRa4lo1KT4/ASkUNlg2dS6j0VfMlfVbMt4gvEDjB/zRHNUORM
T14OVTtIzoS/gNjrht0MCcz+cKjrtkY9LMsJeQeTsUsZ00y7xMb+Gg==
//pragma protect end_key_block
//pragma protect digest_block
TsaFPgySySED8DOfkJpp+oTO140=
//pragma protect end_digest_block
//pragma protect data_block
+LHzPOhBXkcdW/Pt7vmKPqat1GNeScR9Rdf+I4weVprMToYAzf5i4UBXv2ijfBGO
2vKD1OTeDMnQJhH1CdPBcyCWwMHp7yxGlz1noDMOSxsk5Sj61TlD9jFGh08sHm0j
WL5VqnQlXSFeAzivvyT7+AFpTbGuBffebUD09Xi6TzF1nTPFMxbd3/BGMgNolXHI
q9EsJuB0CGZ9vkK47BGlkqY1c63RkVGzCB3AoajkS3VLWlPu/8jFclXfg47W0rXj
kkVXJqp/MBOdRSZugTnOBYDPWsZlcWQeU1K7xggjNI+UKSfWO1Fv5ycJmnPeJPzO
Y+bm7j/7dVIcOZpNWCVJLT8QLJlUQ4HC+OkTudiDZMmmTFxu1Uf0djdwfaTAOAeY
Fpq/ehlcVP52XT+FnamV0Jd6KDf/BQ/pngWWWpyGH6YtWm1eWjo3D8ARtmjodEtJ
XlSGjnNY6rkn3MST1HfjQZancAPLqBY+kKqfgleHYBzv1GcrcssvzMuZLf7+WxBH
tnkTe3DiarM92tUmToGgZkz5AFhb89+1wr5ieBgk/wdAJu14de/5S68QsZDXr4em
b0mF5f9HNwaaXdVy3V3ATTXXSfTS1m5kpjSn3DPKK6XyjNx4+r1UXExeY2Iy5Fhd
xzENv/udX5ShJxxy0r0QO8YW64YOCpbk/QbztgsJQpDnYOXh244X7z4cZEpCVJgM
8U2Vt8p/XZQCZQhaQf4ULkf26tfdY7o8dQRKviMNPZX3L60dqqqbw+tzalav/ISy
pe2wt475GnqMiRTLE/Zd4J6ELRO7pTd0GWTegf5h+PeppOsAKuj9fEWOUG4IzE0l
Na8r2iMJH9+a6uOseFxgCVwi347t/YzvTgJePhKhIQYHp6U6naPrk8ASjI8syjvI
yfLGvMNosZYl90XFX/xSKu3eJzYsACL8nbwFG43Dkkv2xIsbcyEUOKYPgyALgDta
yPzOAS29JOfOmSXFNjRxm3yAUa9IQcDjp6qyhmktuG2wNsgD3rFpPyWFepGdLxUV
0SAAkiCfMCDZIaED1gfohOoqBC1dA1C7R428beu4cSLwyqWUYy8l3JNMZZo2BmLL
SD0XBKcv8pE5iS72/WsvYmUjGo9Lp10sP8qlagE+QBQBvR0Oh3bfJpChfcYO7P7H
qky+6srFK9UDw5raF3D7dXN6BfN4IMTqqL4y3ckXPwrep7KPW4tUiAfMKtNojF3W
le9VQ1vgrNXBflopwEEIQ2PGae+IYv4nYoTjXjMHXmiMKHKHOTluv3imPAdPuXqu
8nDVjF9N08lQdy9d2aNWTOSYi6wrloD/rEek2sWXc7unWI7pz+Rk7EL+rjbPCYpU
lLw9xLD/6gUz1zNMroSRPZsv9SsuQ5t+MzwWaO2iuQslvOm5/ALy1GSMwuxnlZJQ
nBGMgUcspvmwH54Cft3Fsi68UGaxKt2WaCTi66v1e+tToYu9O+o13EVXwkr9kF6E
WXptSwhS4arXJzoXupVodigKhQhxlZcEg5nliT9WUh7P1xJaU5plKhoEA1s59vEO
pV27WZsE75Cfs/VT2TV059ZUS8LQMXVMTHK62QCYd2a9lwWw/UsE44Lcs4EHLC0m
CyUiGEaJF7vq7ECU7slQ8OTGBIe69cSVKc/wVx56IEqob7Obt+y9zwvfPbHRxREh
z/pcbvEqgRrz1EXUN9HZXY34JKMKHaK05Qi+hdmBnNmVhQuzMca+Azdd4rD8JuDy
EGN8mX9k7bTKESpcsQaU71UO40Qju2ftWrYylx6gBDiIBlSgG4kVHsO6cIOFuf0/
ujf8o+WEdM9xsm7N71ForU0211OEXfmXRYBVQTMJKK7vGQqMR6K/qQXwFpX29FWT
iI50EQjz/cHeUN5SVy+DNpJK1SIKXAX7yKTlluSNmrqvVHdFPdai9A8PwomlnKHB
xqs0tEa4EIqapi9iUprU1qsMLLVqiXwtzf3v4d7CeR2E6QrKmG0GdGIYM199TZIp
PiR6c7Fqi/hYRnnH0R/z/4VIav6QMdZ7Qpzvl5EuTINYo01/JipGmDzRpxSg5JAA
ikpoHlO6KqDwrdzqx9Xt4Rue0Yyt+mkSqgxQykYWrYsR0DCwZkfZkuzrvwvUhDMF
VGZ/cDWJxrt/bxnudLxRXucmI4bE5hU9gf2STQEOeoE+fL9ZrfdpW9WAJ/xGcwJE
cfpuxZHjx9buo03ToLYUgs/KaR75BcS4KHovALlet++KUjSLoWzDVdaqj8fs3R7b
9kyYD9EiMV386sCfFBUN9fTd+iAHlZHh5EMcPq7B6ESVEyVYS1GV2M34hJTPYpVN
zSFfab2u8UBgxETOIFs/J1vyxUM4LK6P11LcdRM5nhtZGWmBLaNGvR/X1NsjYBm8
vSgs0SOYDomG0A1zlAxZ4rcv1ev7SKfWGD3FXT1nxrm1PwX5FG2qafc9pKsAnhXz
HSvDgz1UkFfjjHEpG9GNvL24DzffhpF1vXAFbvHaS8HXCFIRsuHNqMweMFjS5tDi
XvFkiVVxqhceYVtRU0duyjeFxhJEIXudg/Xvi2iFjo0075hCduzwBd+qbaXAqUqx
UgafWPaXPatQ0jsENh0Jg2q2UTX1lIgS0w7P+ioRVHRLl3ua8rdlSn7fwhtMwXrU
L8X04sLzrEWH9EnsKkdjttMEapF+JUbGfAJ1JBcGF0Eo7/4HEa2Rx5u3CeegKgiE
KbpSavoMBWUrHD7/y+vGNntI8o3yGyk43RsZ7Ua+Uv8iqQlEPI4OHlj+Fz2lzozW
FsmA6qTq8cJwjGho/0wzT7qAarghbaqwTAZKHFt3awBGgB4aw+Ur9/OlY8hj/ltq
WXeWEHVeaOcYckCf4N7vqkGihXOiq4wPjvOxZv2+XPpsAHJhB1/RaLCEFVFVuu3t
f1F/VB7pSU5LW8wqb7jve+Cp1kWP3ucvR0NJO2YA0Ay2xsb6PEHft1z/yyoMDxOp
rDgU6DvRxCHkDFP38akRc0ufIOtq+W+686X/3+CBUHhxDnOq9b3qqET3u0GJ+jF4
ZYo+VKoJXRluM6ofFm0hqAqi+2KkZGwvQzygaFYaVWjq1z/6IQzIJxwIiw60lkcs
0e0et07GtAnb4MBgwIE62xdXOGe9bEUqGHiVwoRyzfPWE0fuVfMVr/3pbSR9oUU4
aj+FjlwRRyOm/EqzRGZU98mjrqNpdXGKw7XASIaITCq6UOs5l9xUhchjqGLYjYn6
c+61oFacLpEiegeE73C8aeLRe1xkNRJ1QkgxxNHtOSNxH5wZdUzUDkf2W7w0335K
5YDoptZov7aSS6J7NlNRNLxfF9e4f3/JL3u6cAfvyzx5h7QGJbjGdrdGlrSn8YuY
EZPsSGdxg3NIX0c1fvZAOWKCRByKb24d4NA8we9udtu4VILFqX4SRR1b1M/voZtF
r3KLE+wWaFcfg7lm/TL+1vYTm98+L2NPgkuihVc/YWDqC1dWpprI421vqtfmEZ4c
pgXL9hjQ1bfy4PGWBrGvoIEV35/W71vJsPFg3TTMc7SWaEl6xLzRwkIVaOOz45RD
3WJNU3XkCWWb9N9zKMe7t2byjXtVIoQrsjVAGxEHOVvapMnEbUFiblla925BA/YV
taqWU/FgwJl5DY2j76WLDNyj/PTXNtclNj+sSCTX3qPJWNb3OCQiFySoeT3RJlV2
BIFPXzGnNzAxiLv117/RvjY6SLeX6ahFnXoWMYcvJvEW1rbF9VfTIi9oKn6doHHH
DhoI/cQr+2xIJ3+/Sgv95ue4dB+ww0iEd9VlZ0kt3k/5fLqz1Sfjeaw3HMENCbvn
b+fIHtboCTMcG9k+0OQ8Pc3hXwfaHX/yy6Yiyjz8VLVASQewxoetfY3JAXAjOmTY
K6u3kEl3V/jY8qsqW7mwbCCKS7u7YRZo/hHev9MRS+775kC/h3R9mIqKHrZRwjyQ
uGJb7Id/+yZJ4kWAAptdtuTT1+z8Cbzv63sP4LxKR/uU+Gn17T9N9L7cmAKL/Cvt
HrHy4zqTAWAYxlJUaS1EwXrU2+ofE4Ujx5qMwukPeZj9WSMKjR09nwODyjBnD3dc
zXHHPPfN/q7gr3UJeGM0vxDlB9ttLY7wDyz3iV+gOTMQqeKKT6JGmCiMwr0ic3DF
rAXEYTnhr3Y0lLzEoX4Zvgb4vU8GQvzYjcnojkZHFPuV1biS27BQyOu6gvubnN3L
kTnTA4RKNW9i8WBLc3bRWlmQ+w/3R80uD0c8PgDO6vc2u7bPfqkbOgmlk+jAnt+b
4Pk5bc9Ss5jmukLczC23231zJv35MNFQgmQ5LHK07Y40LxXF1o394bImuAWhNWNh
mHwy1tJsmZfeqem9XbAFAZU9UJ05GrY5tiGk2blsOalpr84tGMQJY7B8sVQ462A3
GrvL1ViBNvreQnMi6LJt+km/z1gS6IVulgW3Ghwo4kwc1z3W41U5NQnOI1kN4a6e
id4Z5saZlI8Z+SbV0gB3WL8g7UFkhawUNSaKpB/+H8l7Ue4nYXOVPrJ5yVJwgJly
QaHwOZtgxfq24K33W4+T6yKpvNoag5f6FhDQ7cITYGpJINgWU/B1Wr3cM1pXmkRJ
f0aOiC9I+WYTf2lryceABqqMzHqhXuDleXgRDCR/TE0KEWRH6ZtG6jNlP0jj1BHi
p2D3ci77YdeXgFhkoW5hXn4ZPHV9J3Q1Ou2S7my2FcizK2Ljzzz6HLVceHV0jkzE
5JHDBg7OngIjX/KD5+jJWb+/JyFi4gaxXTsvBDEgVmZRhjDrj0xDgETr4MoNBLIv
2VQ7mEAYaJgn4XyXCt72qWzkDU6neyl30CQL+PCFtsPEONYfa8VzxkomaGf8JRjl
d6j1ZzLe6QtkFVHxwCksS3ZkBZP5/KzWzhi2XkW/eewt0C/44FZi+b+rIhCgqf/G
5U+SUXsE6wTbWbwyE5plmkAjqoWiAWh+jlor2aA2QdlpRN070QPHn2HcL2R+ufAq
TDHt57MfD8JdTPF2jTpwb/Wf7Y4bzWbkpDUK9R4QDbEyF4v1CoH/PFr3efxw5S6j
ot3nHm7nh8xfgzMQwt1a9fONQeFRO4ybRgBVnKhPVnWkNwZwhOQqyadiiqzaiRS3
s7pJ2b8KkLk3DBqVIyu+fx9bQ4GTubouNgqE5m8V7pPsUiBKpJ6iJxCNQxYBgOE2
9YZJ3KtgHmrq5Wq/fmqnlg7zLkr6oZTi6utyo3xuZNbWhKMRL8128zKcMBSPh2c3
jRixSA3kaOwFvXvtlk1FQv97LbCwBPxO8CCYLf6Zl3huMoPJKnGST2oenm+EHcDW
4IE72/7g9ctvGfLeSoksmocJofmMMMkJB8wnMUJlN40fb7jVELSgabuSXDshVcyq
Fl7uwWWJ24l/dmP62cnkYvU4sV0y8hwfurHwrxmhekTggbHe2A4RT2IR0NB02axy
nqRDUSUVnvW8Wje7cxHMAIwqezSFt4QR+vH8wb4LSSIgbCoD16G5XIz1NuUuVyzr
nTb1GiNvI2yHLX0rW2CqbSvv/CKwx6InngJZm408C2NFqgvwYKUy66LGug6f0xLT
lOp98QAVhNYRkX3tDn1j3MkxcoZtzG3e9hG7HSCgeXmz+ECQT1RzFvXHE3GxU/mo
4hnoHBBLFdWZCEPouGwastGZLmpf7MT/N3VJc/TRcYuR8g4XkeRc8kzonh9I/QBi
DDQObhAy2PfYfjf1TjFCHdmTeVgL7KzAamAu42GUrHWEo2tZdofduNOu2TMX7sDs
nopMM9Hmp+7qGUzIOsXEAyiMZ3y1MP9nn4x6gtaSgoabW8S7WAVVmruvvf6UQTck
Xkt45x6WSxqA6odnFRG8OEyuS+GXXpWSRiBEuejkw3DzXYb89tp3v+tA2fR+EodT
rxf9MyYaN6rTlJuVFjFHwl7G/sguZMLNGpdcE17hAGylzu1VbQoIzKSyzk1+kmzS
mVD8SZyg/SIWPFK+lefgegIUiGKFSYaDfbzLbvfkxADrUBzPTEsZ8MLqqUqdehg9
FaRgfz2wioA9FKpf7v6qoQw1XUdYEXW8sOB4pOpab0+EqPJPBl21vrqdmSdUK1dr
KnUji+6qlZ/41lZ6axMgXjWkOGTAKXT8+4+BOdSrjaRSQrnqn57tkv3WozH7oc1S
EcFCCQ1tcqQI0YlPKa69RTsd7tqOha9Z7UJyuZBlCGeNnFgMuz4yKUPneshH2Oeh
nVCawRfDeRwTnr7CXHRH27FnTzj8qabbaRwbOc4nOuldd/XgN/9yzAO7T+Ksv1us
GQ0t+8PT5nyqJd5dom6gGIFwFuZq+6Cw9xWfGQjoZ6t6DjE6p+PGO52BrHuSRxpu
MBIc6fICDo775myoj1Bimdac1zKdxKWGwGARY7c+kPbxHIgVVwET5QRPEGrHe3Er
6G+AuIT9E9OsuGxwMbdhrxbPDEA+vSEh1ZrTs0not40ektScy/BOPreuEHT2Iqcj
KrkQ+lrljukK3EyhzmFfszCRzoB5FlPGMc4nuGIicvY+X2SFPlLeC8p6/c1bHKy/
PF577VEo3AoQMcjTlMpdEEJM74PaIjme4n7U3eb2T5yjbq/hrQ32KU01BzSLTMdK
J9W1Ored8gOt8Gp4LeJM4ZxGXWkYEcfwXkcoh4fUOe3a0lxbpJ6ua/JeJowXxStq
ggwFFeqaR9GxtBlii3oW0PjkqYfyz3/gpe3cqxtNLZ8FXfNkyO7T9VH8JMgoaMtd
Q7geN3mLJ0aHeayT8wGl6eR/6nU0jmQEmrBO6f9HDE1pOY4QsikkX3tIUAu1lDJN
2wdap+uvY/R/D24ihHpSvEgQwoNMpdTKvqIjr3JREGSsAwV0J4gb62W28hh4JTga
gCn8GRoVvTbcKsiVlY/TIeFAemtkC1R6du57jqwOPkV50f8oGTyoJMw0tO9YH3Nx
kKMvDkfolSjSUOxbwwwN/9FpsCfztoYxDOnNzoL5UxatjOYhKv2v68tRvM8go7Gq
x+Se6QQV0ezLiqKE21lGTVQ0rZs0BmpL/e212eVEbc9QvUjRkLiO6dinY+dQIhFd
3CJ1lki7bzEO0K3WgH2AKIlypfNs3xqjfQUj90sUOuEuAqKSE+sdKGnLEfYLJAWC
8QFyFlt00pWiuuRGeuVTDm4PRgXjjxUyIKKQP13zhU/vKzUseV2Inh4e5DfOq3BW
TB7XQinCH5xUexyenVgHDZgOSPcuYUJmUs4QuBPWZtF0n0Gzxtv9WEPhd+zOWSTr
hVQ0z2pqWbl5bvLhRvqxJAco8F2eqWdlbGJUVuT0iwaBffl/9q4rsSazs6ZIYQiP
PcLZaleosjWITK51RHTk0wNJFZgZtDhEid3WepV7MEyQo6xzgJPR+5NP0knZUB+m
bJHN+ZOClsJ5LpiazpsESjDcd07AiOfmF42hAwJl99x3yq7e2dSn6XlycR+tw2Yw
bpfJRoVFNcbrAW/6JuVzXUvj4k3ryRZe2T7jzcAPGkjFuPNf3+iEFieiU+9eclte
NGWdk+efeidGFxBhlkMYBB0P0O+1VEkHKjs5IpkxVmENR4K46PUelDR5ttS45XTR
yYJrPrW9wfxJl/VXxhTPbeNve1a34az8J59D0eZP519Ktbl/99D1j3Loq1W6KDBL
7+YpRG5Fm+RkJ3dIw2KsJ1tIDviNUXsjWICdHlQyLveM46MqZBlyt5WPucDQ1IPL

//pragma protect end_data_block
//pragma protect digest_block
e47eXs9zG92f142YM9jflohNMx8=
//pragma protect end_digest_block
//pragma protect end_protected
