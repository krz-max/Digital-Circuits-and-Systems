`define CYCLE_TIME 10.0

module PATTERN(
  // Input signals
	in_num0,
	in_num1,
	in_num2,
	in_num3,
  // Output signals
	out_num0,
	out_num1
);
//---------------------------------------------------------------------
//   PORT DECLARATION
//---------------------------------------------------------------------
output logic [3:0] in_num0, in_num1, in_num2, in_num3;
input [4:0] out_num0, out_num1;

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Cavv+/HUPlWR0l9dzn7xZp6AqasuLBLtZrRFcOjlJ9uVi0MTIVdAszUNPukbJIm9
e+16HKb8bC6ljrqJ57Nj0S0PSE4zjUNxLzHftacMn1fD+JZ5m57+mhQxPAnO3Iob
H3ZDsa5ZIeqUvQFLZDg4cH2PdwikFYBXFRWLhkp/GQMOYeB0BQM4Wg==
//pragma protect end_key_block
//pragma protect digest_block
FeIJeKhc0uXXWf54kZt02SLWRXQ=
//pragma protect end_digest_block
//pragma protect data_block
yHLHsVitzUzDWXKRZTSMZMwLYR2nHzJ6Qv5cfkrtEu0zwwA6hPF3iVv/0CvpqZbt
1bVXpfQe1dfeZVNw970OHoGsIL1yMuALpzmn7tLyPmRAEgTqlMUtb2A2gwtyWfKA
x+CfUclOo/iYF365iFVEFYoooE+nVRB3VI+T0LKVfM3jzCyUXI7gThR0bUPI5oYw
Ah/AnC4VdEjNzaHEjPSmG+n924aMt1SNUtPKWNAcutuTfnLAOkUAs5Inig7erYnj
Qz2vzsn2eajoYXnJSz6YtPY8QLVxTVKNT5+rIjs4wS5CBaR1fDdBnAwBT4ZQsvzx
uHOGWswSD+XHCVLpuVilP1Cqcvb3mU7xUaiWvU0006KYxXQBk1cuiuKiHpxYBhRG
VEpHAiwszzijrxG1vlB52EMBWAwM4RZvdTcCT++P9AAeb677g5B7wDHJAKw/LXZb
bBCtus84OZKGW0x6VJvlswecPjH63jkHB1L/u/IFkW6NessvrM4aMLEASlmMxuPP
jGKNM0u51B6u1nKULewhBu5cGsxDdYvrL3PMGxpT1WYAKR57PKigY6K1KJ76Zne3
2+yA8TdmhjIeyUsmGZU0MOkwhcMYM1pi1ak2lUUYtX7ulMNYa6FAdhGWeH+cCVwe
Hm4CT2ARInC9jXLxL07J0R9PsCGf7uSYI0MCqpgHfP27Ycp9TOT7RqQ7UHdPR2g/
eHERqgEnBjCR/hkc/n37YCcyJAKvXfrjm5MQRuBtJcRQkHDqvHc7/ekgml/5PMph
L7g6TSpfsqZb3O35Yh3HOuABrh66C7j0GbU5mKk5Hy6Dxz1BdQaep0pDtcRcd2Fp
jLZfQYySQmx9p47Sd8YeEFeS5x8bCkBrY8YY+cMZrBMoBmCRkl6CqZnbfus2/baz
Wc14tWvLs6kVcaqnaR3y/Msv07wYMlGAEHQRNI4QicAKArMdNGaN1I0XdEoCduqv
kC4doxX1W8wG3gb3eGEwFScLktWaDJOj+sHYfwZi9RmavcN4eQNH4U09RMhzbnsk
Jl8CCs056peWUupMmlcVoUob2GgOKHJyLCIIYNH50KPvvVMWZcH9w1fYRRNlSTFC
TbqO4ChNhiydSlJfwmtpgXhmIPd0W8vpzol8Q3Px3OIJTQfuR7y6+JE/79/4S1cJ
2LakA9VNIEydy6srYyaCB6zAH57EDdEBMQRje1dZnciULiv9cLNjnBJSTFvA5clt
JlHo2Yqw8wS5O+X9O5PqF3r//YDdnCmgg1hqnE6WyCb9m4OdWjlMTlWrrRwMhpUw
og6soho1OHzZwZwaxBClz6f1hZ0ThaNXGmVPhBKZ2Ml8jGmlnQY+vVeYF8ercVuT
mbacQeS/M48wsSF4HQu5SbUOaSjYIpU11xqtwxJLPe4qeumAo7uunP76y7sBSuma
iIZeCHZvgR8ewAjUMXY56/wG+vIiQACGu+J3nGnAMoZ3dSAReZr8k6cOY3/tE8JG
vB1xhV0Wizuq2IsY6esTE8VecLmJZb6y+fsYxFiyteO8USb1z8449RuXbovzf/N9
6O/oTBe5DyFWyj8gzlxzhyUNH+8Yez0EwqE3FUP5QgR23CWiHLRUlP3z0RA8wZTi
aOQfpFYaeXx76itHFdfze1AstA0jQopF5IVNX7O7qyRKL3LXCL5AVsFThJ6G0RXU
NDXvAXrW8xSGxPpFP3jA1ymKpfmx16YymPJGqif0LKftZYyTHFLnZbatof0NvHZd
GrODoBZE65UbxhjuGpPNCaukafkWW5MXO4zPK1UUud+aWEpiJKPCD/5JzSqi3fGW
GCDmKBbL26605yFletIy+twofnzPhuafxRe50GkGJVlHFg71na9DCx3PJqW9zSEx
NN5Jrf9guEjFks0dFuTGQyHUQYsM+1EadAhCFpxI8FOuZoSJEPwKH6Nwd4k/wMP0
6CLUONhQuwlkPhcQJTTPH2uP6qRkfMpkx0kadjWG/GFXWOzL3ZW3eYrAEofl6ZBU
gp0FZ+yv/c5SU/CoQkqfxp95VDYIyG9k+MFTVBOV4IMsx9SoKjrN+HyW4QWUzNXW
gyHXNVic+BSkAdlpROy8Z0chBe0ssy13cz60LaL3rua+OhTUz4kS01UPMSNDvxfr
Q/Bjdi2YfYtur2vmj7/A6Co7jmw0V2dk3MJLXy7ACsmvfZAxks5S5iaxguOFTI4m
CnrSmRnZpbLqVeGp1SY/MLtZ8PIzTwgSlOmDtXyWxGBc9aeMOEUHy8zRJt/adCLw
5gV4kNlO0QqnwKavP7ASTTYQxQATGt9IJ8KWpz802vx1ti88FzZuzTT5tKN/3mbm
tdo0ZtXbrQfxKesQB2YRckXQXt1h5P9qEdgs/NivQ8L8kLCaHziJYdjBp8kj6YfB
+51j8yTQ4hZNp1mzuRiQ1vsLQ8cEvOxWhoEI9P9XKLaVMMbik7TYuqC0DCJy43Y1
0LMtbN1ifpm6TVaFpWA1j+dbcVRSd6O2NCzbfPTI4vQzLWS219TL6c/z7G5BkIM4
36AMwkZSAFbcLYHRG3qDnAZhD4wCDZmJv9Ol3ij8u6S4gwwqDX5hsohSXCLgMfMf
Yp3xybRqYrvVLcaXKidQp+uB9RqEq7cncoCj/00ITKiSl080aQVjfSoIdlwsRZbF
TnS5C6YqxI7+hDZH7xNGXGZjILUAk4tCC+7ADEnY+mVzRjgad6XoTZ+Um21C0lbp
kCNrwbLIfqdxAZQ/IaV0vvvD7JAnC6XuceJiv2OD7UJUuxUldvedGgduZzG+uQXU
/HZDTFK6Nk/mlqrK0tI2byYhqSQeewHajZn0JC3wEjzP0PrOGubtrhdZuK2Xxdkf
+ed6RxRJ9qWIFEPtfi91uBZKpMSJqi79ZDXO4iU3Pa31YK/yqwU0UFM8w1BHvAov
ql/Bz93J+FrvFMmqLmyxOMTvdMg6TgjffD7e1UK5hV1VFSsYTSXs9InpbNqGr8nk
JjFb8npf5fh341FHCLc8StaQx0UzKRvcr1Tgk0cuKDtztL18KipYuXVLd0Ab0dpI
anqkHWHNJceW5hkEHgxG7vhELtYnZLE4er6ie0acSGZxhl6k8qZsGHt7qUUBp7sZ
rT1TwJdveAvILKf1WQMwRLaEfESDHuC/1DngoYWhQEL9GePQgbGh7r82pzzeTIPG
gMuNjZ19L0VL8KIZwJOlqsyjW4tQV68jnk4j/9pK0G9gbKchLHdXMuRR+lwIuBDN
TedIl+YS4QhJQk9HUjve+LuQJTOOLo3k/Vz4cX8ilP/8K6obnbpBS2qzX+KUuFpr
wkL3dH1zb1XeX50Kt25RBzja3NZq9VPkIjch23o69zveOv/zHWRnHEL7+8GeoH2P
f/cPa0Mco7Wc63BEbivl5Aw2clhneSu0UYo4Pzx67jQjKCgt5oHndNx/2FuIbNe0
PI8f0kCJ+RpX3BP/Uunku7x322vJ90CwzVyB0K8Mat//bfU3tUwFt1HJxFsdwncj
x+SOvePG7U082BLtSQyfp0DyCMXJYchhpTSC/vc8yahbeDUwFjSNJsULur8MpjFf
pnq/BqsE7YJvrPoObfZQnR7v2H3xq62wDRHoWnKjzUUcgkaT9+AJ13F33ZK6zrbl
lfKLr/blxOl17nv9PYhT0Bx5Jq6P98jIYYiD4WI/fUi5pMUQLfh7guz3ws1ZmKxe
ciuiUI1fFRspEZ2aiv5lrZkNSmd1BQnUMU8IzvYuFHEoTHucK3LcwZ8Au4EIeGw1
MQ+uPa0+rX6OwcmeTiipLyBo2kicjRRPUqrBXCb4obw9Az7wYAj+T8DCEOOrMQA0
x20rxBTVT2TwbOODnayd4TQNXzF1NhZpWppzLm0nQPJqDNQY7gj06jkym3So8jYu
8gttcf8EikzuxMd7IaI0s+rOSGZwmKMrKEqL6T35rylEsMRdWe0tsGtHEXGWCXgS
kyv8uMFqhyiQMZBxRw59b0CO1wAN2D/XR8uFh7UdvX88X9QzofWqyf+KIsORPXkS
LbwdMPr7Ma+b5Q1mjNE4Rx1gkTFCHfW9A/Zp76jDR0BwHPkolgIJFE5G+VUo6+Di
2nGSgpplN+BN+ZdPm31ou0e7YyzX0ghUtaq/hZu2LGSOpgeKsIg5gd+J4FI8jdDO
lnq+dLC0ky84QaTVJtuOXsIQDTkWrpyuouqObTCGXa4smmqv3qtBd45Y84s8vLU3
bSbNqS4M0V85RZ8Rs7JjqtP1ay37VgNbQXzfxxo0tT/ywyr5vwZA96tRzxnStf68
+jvpsV6NsVr/79WlYOGddgw26MkQZH1wR1ma4oQ5LJRcjTlQ8o2IGTd8PSTdyo36
oc5CiYDSSdAkcMI63nM2js984v+9g/yQ/VcZxKIApw3ORFVu+S7TU6UkLT9sw/oT
vGapkViNJkFRCPWeohtmTHYVSiqmEVfJtE42frBzQDVam0Q+20ijPdp5HN5TnJ8l
M+i3hhw8T0eBWZrJZPef0JXDu6i/lqRcYbMTr2hQTyBYgoUHEmSSyChn6LCRV0Zu
kgvRCAx6ix85pgNY9QMvp1aJr/j4UbuLJlhk1eKorvRK5WrQwCZ9W3XiJUrKfvaE
nV0UvFdawcwKItlRYXO3bSbY6ivPOkTE1FOqxiTWKsKU9k0pzqd4aBQs50Z2E68S
gx8AU7tG57wNzsJxG45Xms6GUw0It9LffLtcBA8/Oc03DFt+glphNLAREsuEmKzr
Uva+Q1dffvyVeW5wLFcRBDIrcSH8iaDT9qMctF7aNqbqs7W36lyDfn84Gdi4LzFf
a9wD1oNAvE2FF1zvl7YZwQFUff1LTb1T7t9bffMgeIpZGVrQxEIbnc5CrGRPZYxe
KMfXSQHimFWEY5G+UIZmUyN7P8xEErAr1FU1JpJohXC3L4qhKYbTHjcZysYOuCoh
Rm8oaDcCbAB9x1YjVCg0j9ddiX3DdqAycqeUW8R7/Z6GsyO+zBtYvmn+n71My2/g
EqjmB+x4XD0ftg76isD4wegeV2xcHenJmVLQ05iW4ZtZc2Qu5UVDbLz0+NsWT8Tu
uF0svVxuULDUpwoMgPRMC0E7aY9tJMEZcLx620/fKX6SrhIi9pj9PWVA2VwnAvBm
MuDIT+YKZ+0pqhvjCG4C6o1qwoK1vzu0PMWieiR/3AfFXar0sSgYXRKZkpn/YxW4
r6Jz64KL6ZJxe00/9J0Z0TUb862hoh6YL5YpCIsvfa+VAFwuppsusHwdsNLvAjWK
rb9nPiTxecT1dOh1wjg0eVaxB2Vkw3TOJCfCDwbxW6HhS3NHZKBuabxZv41zr7JD
kEoTHyrKcAwS46yKnnvrku7637V535SN0dvXnHmxDVj/jFxwnKwqNF+IDXgYx08N
swOYM6w723pV7pIM+8GLxhS9J3cC0IckZRIsPiAMg5vx26Hw6Sfpv42MEzrx/V1y
8iWdqP5B3XL9YiFPvJqH7wzrl9VEOMVXmJSSXeC2njAsjX30iLMkAK/aV8BzfXsN
D9DYIOAIxY2BkL+gpu3Qo6EVHTbooRvtQuk1DFpgIUKV5qIoshHwC7QHoPK3RpnY
9i55Cc2x0dsXEgs+SEH7K3AJITBBy5RwOsohEBy0Mjdacu2A4YbhLAtSxdd2X1a4
sHkukxK2rYR+NW66jpx1RkiuMLULYhxzCQ+nBeoSI39LizC+5S13Tbu3lr5bq+0z
yEzWMmGCNxQB10GZNNrHjBAG/nNJLvHbv5We9Uj+0fkYyNp2hf4s1+E7otHmDS0G
fkqk4iljTePE4zOPx3PP8ksYFRy5vNnyiI2xA3yfa5IipAc/j8XPXF7TS/psOREX
0myoqIPA+zarURkIra8ZZsgtIL9ecrlY5iV7cl51wsqvjEgK8xvOq6kGey4Xp0YZ
ZXFNDwSJR9TBX+KSf01Gn2J5EyhSB0gFhs9l21qv+JGN19/yjxjTobafmxWRNNt8
6mjub4xeLT4YmB5CqDArb90tSLjgdEiWPa3vhp7OYy7KsG7r5frZeRxnAG7PpvTq
A9FM9j1RhZQT8BMSw57fxui9DGhTx5UaclgFjB2k65FQqb6Ue2/FMdwcLVN8Sd9N
nQnl2Zgduq6uko/83aur3e67NYcolmz1pC0aKQaHEnnWfkMVqHBxl5EblrVRJ8Lj
pixQu5lSyQx4Q3TpFN5ePb24GVsu0kH5HBIQI9yJwvRz9Isofk4E7zuasaaE2i50
hfwqs0v23Xllg8Uye3mPYXl0yue59byQvKxEZzCc6AEuV7YrTkBCMmrA6Iqws/dT
wViOtkGmRai0WjKj8mGGrkKH+luCcM5i2ukjPc04N5uhNdau8rtNG3Ga/9MUnVPa
ikHqVrBVMs00ELM0yTk6u+pLCs2erWqNDKIRFHTo7gadRCVd7hDr0FnxWh3PgKzu
oJBsiOFgQs+YCsSj5CEw5bEr4Z9c+L3Lc01k49VtUGFRJTbS/VPnumf4WMhmfqpu
0E9jJ950vkecagUTGM/0cSX4BIUZBI8Op5XI//OwNj95Gu2ppFcTH3qgNApPGUJB
yuPgkmA9htkvmpirL7+P4xZbogVJycy10chMfP8Q9MNjqKtSjE8kPwGw0MOKXk3+
4wxzJOPSQlKqXAOSgkqvpfWnmR1Cm7uGJdVsDscZRJcS/h8EdpVzmRRLsGn3GcIi
O8ViCVojTgh4qevdKc7A3BfSZzP/2T3WFpHd7wvEWkmTbI/x4OVDs1w4TjY2xp5J
lDcSSk14eOwKwk89gJHRtoZp1xemtTQHMlo69yhzM6zN0wpri1nnzy6tldAvoz21
EiKHA3aOWIUt+9th3dHDHwijV9jyfcWvReIXuvRY14DcARRRgsbRSVFLZ73avVUn
OGoEJuTzjgtKLjwMtq7pTk9qy0LeDmZ4vqhBfwwYJnRX73m3ZhlaqGv6/vuZ62aY
jCg2b6o0AaaUARtlDrI5pyc6ogWeaJqibcUP6Zr76qXttBULofrWgOsVp9l60Wvi
dUReaYwdiRzgKOx7FLxq8OYbiHXD5LbF8Gcuf/tpCEKnZylb+Kc68Cbisd9UJwUu
bEpJcsbV2Pr9CXb/jaZ+w+Bvs1SvVR1jW+2KnhoNC3B3L3zlRV5S7tEChO/FKdzI
u2ySzMm5xBpOwZs5I3Q6fP04x1jiSoV2BJo9T+pbLLWlaA9vVCkvoTJEG82z40ZY
nItE554yKIOnaS8aZ1L1a8HkS/mK11fnXkcj5JCrCD0GEmC8r76PwA9Yrz+CaEKR
3LNAc2iozqaueF679RNKHRTyVnS2pwtleFBG6kypowqRrogIt33vqdPKnV7yMOxE
t6AkbMsXfuaVyszMXxUHocJBdjfHS/u1empSaOtt1J8Q70bK+6e6c//EiKKYo2df
1wm+lOIlf0bmD6ElQwEhZYwZBNeRoFIXhKscB0jpRQi5KMvqGcWdz7UKBNfnLW1Y
9bux1Oa+6wlGJzdlBK364DpaCtITBn79h3IeJiwdi810fv0gMn0pl3WmEvOnBxzM
oGPm5EBt6Ws6u2zIYpe/qm9OADKdC6NUPRM51OlpuoGtrWQaGzYUNXczmRXDzlxY
3SQeGV5ndd6ITi/0xpr3YLCSJwSPHVt9YvLM7RBtvS/m8lFZIkBTysKY4tzSgxv6
SRBkjmihLnXYqQkGjAV9eshE2bfLita3OpLJoydAd8Lt4KG1J95IlvRFBsFp7KHK
16dfj6saxNQYf1MqJgeQpiESAYZNwwM9Noui7/zNdN53HynXHBpKW4RjjwJOUAHg
AgcrGhnfW01ymegRM2AT6g0oz50M0Zr79G1rkAj6A21NqL87umEbatDAgpijjEqx
MYZvahg6CJCkP6iIhzVaWZCAAI36t6fUCQPFIFxV3DS3rK4bbJaQa2g+cyFl9M3L
EokdE6Qk6eYwqbgwaKzeQR0SMpqR5E44kqFX0eDouXC6RoLnMbM4hMtUhSpY7PXE
SWJyQawSUkVIZFF+vQaNeKgiR6ak0DRnX5Utb6MqqLlBFEu2RUP7jHjP8GHzVZkb
KDPI2cYQnPGH/KF+LwNGzMomvqyz/zBKZzfKmhRgc9ZSb8N/isOrbOaEWX2oBDti
2HsWf/oheXIQZPFj7OlGMa9Xar5FjtBfcvUbGDDazj9FPcO9JFavmXkSYG30ZkIa
UyfX71SIl5vLr86+v3UNPg9YhR1mmDcI7NiW3sD+AUwpiNcdIXjGUH0WMN2Ut2ZJ
koTzoox1amWQq0XxfviMtPHcz9S8ukbA6G94p4SoTd0d99cy8E77De0DnUeBjiJ6
K+BgwRUw7ymKEW8KqHmY/Fr8+6i/e6OChTlSSOr7WYM4LetxBcgxzBrnreK9+yWC
/pHgisnq5Z6CW4TRzG4S4/g60bO4YEO+PWbPod/U/A+lNHIKZ+k9KJYia/Y9oLWi
SQjnls6LHhbYrt6xwJcOcm8PBr6yNKTonGDcmVUeeNaUwKhWbASz4CmikHbm29yH
NFIZHFrlgV5maD/seEJomD4MD5fsk+PJA8N1L6rsWmPLKO+E+dwUeQ73k+hJM25o
zHujtL1Y2SSfyIMLRTSVRR8ARbsS9/X6a3HNwZrw5Ck/4K89S06iq8ekenvofWGS
J8te8kYdXIbWDG0fuPhC+I20EtUlSCRvhcTY9OCUR5ZezbJETgSBzEvdfUpr+mwh
oRlTnKk0D4TF6v8Xq0VGXdA9T+ycLRFxo2WXbTpey+mZ5TP/xwFXzrhq5u27I40R
EkT3m+0iE7vJbuZuVSVqvAdQq7/oSbT3TrmxMa6SMHDb5NlYjF1NfI7aCPGfBawT
NOZ5Sm+WGWhVdsIW2BirhktYo6TbarWc8omIXxa6pjZjFyHjHdqaA4Hm3guqj+qE
+1+hpwYWe5xhHvoAr26CIbCiQYGc4o+z1fFY0brg5ZVjmCGF6rTHC2YPJtUvaaPi
kPvHNBdQW4nPhu87N/HSEQBHoxJRlVs7gIYPIQCI0yEqg4Za0NFjO42aWhAi9p+7
FcUnUqZcxiDM43qD6nvvxt60KDB3KGiniMTCjjoTW3xNohGhrCG6N32Iax/OYngL
vVdp5b1TypQrlUK0zc+vPXK6VF84z5CZVC7LL0Yyd8z9mVem88YzI8979gkalxyW
FCK/Lk/zcBmR50QTGt3/TosESJVKXf1h7BQpcx4zNwOcVTqs+1LVK39zKVTnhEmZ
Q4wdiZwt3OhRXzImfGhuqnrB5LogaZFiZ5n/cPJNwtrJc5ZRFFo6uqQPYqkxRTLu
Qg5CY2D/wPA6u8I31nJ0nGpnDoQdasGdOVBzABFYMhbc6/7sitAUqBdavP7qZeyV
o0OBfehy9DvX+i2tyafY+j6rUpBKxYhUEdTu0qh40FhZQNph65vCWr18EB6Ioikn
Htb7t9iSZxtw6U+zoGJq+3HQ24TDQgCetQja21gpxZWDN2oiM3gWh1JDrg3fuSuo
lpeckjKOoWU4hRu1LS7AMtsQpIs83aPozArDx8tpg8UXHC4x2F9jGU6fkKFaM8ph
MG3Sp4VC3s665KbVaTNfrbl1mXnIcbvDt5D9JIA9wUROrYbU5wvcKjtSCJApOLO1
v95ph0CdZdCnl56QrIxhHTAXXtXbAO941ReIVs/PQsgal3R9zRPSPlaHzefcssKd
PCPi+q0e32uXGviakXk3SUtBWEbCpjCFqeB7cs8ozUzbBNubmteJFgVmpDkIBlK/
WwCatvvhVYtaNcS52zqKTN17ANMW+G9ZQ5uBaWODT9JmZYBCyKYbhX6HT2T02+MH
WkNdMgkV+n/IPgGyg0Orsz1z6edMTOKLfWUN74ffVGz4r1jnOJ75ytXAXyh/GODL
g26iS5YfWnE+ChnRYqCNvH1vbk2qkhJrztFwyxZAybqed5+gTCgy/jWdX4UWG2BI
6fe3PVBfZ3q+InKx7i1CD5CZFOgOPJcjEiaaaqzARvLqOj8o3lhra//O5viv1R4v
hSpNPzbTDxd6YUjdWLyUPlkbw75AH9l+kDMrf+OliU9lun+oQtYtXbRE28knWhO3
fyHFG2Drimttqut/4L6uHJYYO4FYf7zSCr3uJQTiUhb8pgGdcb9x5WsoWpPbDxBK
vEgP52AJgTCL1AfmNfIFD7bcen0rTMsR7DUTfJHbNIJPCXwDZBjxR6FhAm+IR64J
UjDKA1bGAHe3b0JTakCxu40p7phHPyJJGNNp0AQ1g1qbDMHVlBSjSBVJ9bzqfyoS
MyqyvgkogsBd7aXDxIapHcbQNFdzBrY2+K0e2nKhbo5TiaxSHtSwRRW1qIHbUglw
vHev6xoJMZjlL24TG9R//Gnbi3R40GS6vvbs2WGvMsxBE5Q9/M/q8F5o2mX/v5Vf
KWV0/O5i+YUQ68xUHtCIJPgRX5qIzeX7kEoBxqF/2QFOzbxk3717n1F9lajptBaj
iPtk1aCHNGlQ/dWxmXAIGQPV81wiJJu/kSBMxdYQHCWGuyxZ0iAWLBCJQ4NFpk7X
kPEpFS9WGeOU1Snr/RJz19brfvFRhUwKc4PQTKPw43dJi4UGjqpdk47LMdzSw9dc
CFTC1QuAJLxX404ICkrr/D3WTaO0tjUHDp2clGStCjI3nvN3R9uSVo4G4kmDuHYG
Y14ADFBOtDIuOJP02L4MLpuA3+j82wH/PKOOrWmFOE+fqtv3C8GM7uupwH774LbB
09tKeGfoANiE8Any7+TQgleGA73sX8IyYjQv9KsCnLEhYHGfxmziOJrnt64d0c7e
HKF8KIVBbVqn3UdfOzhccIKi+wXsY67e29XG0V9v0+Bh0ov6gK1GHgDOtsmM1kXS
I73C60ZRRZD7F06VwuBB4n5iut94SMhGv4+IdL+brwK5AoMjUFmI1W+74NxDI8fH
2EnswQoOUnkoIG+KBPmYCfuvak0qrptxwWNYcat1AEnACt78k6ToztkizpfE8bXl
BCbCeymL+YXuagVP4lVDDJsdq+vNX44wJD61xKgeHJBxYXRcs8xA8241CCArcrm0
GnfGKWmf7ykRFQGEiBC8PPMarsEMmCHquUBwRmFqq46mLxXTP+HmzPr0+0JEbrF8
TSvgqIqXGHvimH7geUlB/nCLXub2IyUrjomglRxnQ6SlFzPd/IBFWWIqhmu3LBaI
O8yRaT99xOyzRmXqK+06vWM8RWu2qTJa4OlZB1WampEK8fAhCf7WlhDDI3IQ6sHY
xeWEmplswkakCJAxBYPK2PidVgqe1ZlNlNGTpIbln93vHlY9rcf+2iuIc/yi0i7S
iQqt/u05vXDdco8LJ4voPivJnxk4qOFfRbyREPyaWcfNZs9UAIn9otp9DRJxM9kD
sCWJfyx1wH4OhHgQPjqwO21qfp8Xc/TJTPBlOOK6tKZzjL7bTPIfF0PJ18Kcjm4I
TtZe4ybhX2UzRgDXgSUnDRwf2xDOZRgW/m+lnIPJA87tW7qiNY6t2CG4wGP9v80Z
SD4oDLJn8Ttn7h4w8iG1GK1115NRVdqsw6AWIQh78Vnaim8gl6EXdZYSdSyK0473
BGl3f6pVTb0wDRRI0rioPbltSwQ0YZVzVlLwSsiPXEe0QctHnoAPml+b7vh6fDXP
l26Ug5FhhC6L9L3XCdxmTNY5OlAPK7CUOzL34R4388Rj24qdE1J6vc4oR+9jM6Wy
usHGlygJYhSxLr18MGCMnjgaC0voB3aYb9CUs19kSuu1wemHrfoTVdQu4UniBW40
jLqqlYjuyr397RmC2DlhTMe5mXN6MtRR8XpOpuHn452SR03ubmmlMjzUDwPK6am3
D6Tp+9C/w/jotVxloCphHgFYDtR1ay8pN/5nSOV4pE2Gt9TGy+uZiuh7iIwKZK5f
rOwPWhso97BWPqxtIxn3G0ZaCWMYxiJUDPIX3uXLVpJgUOGCylhgFObwg5sv7gHt
yaCblaBycWHlt5hkZI6DtguOSZMDI5d6rmjSeLCp8bpORzhPJ+fsNIusXMTlK7GP
HmxKZ57A7usLpjMo95OFvyokxKyPDwmYRrmCD+MTJzyfIdkmkd7wOIDcVXiGpa2j
m4nYMo6sVAH3qx7QVhGyKXBQjbYQ3AQtVpcuJ4EaF0UHiaYcuTXq1FIoHY1TWhQQ
2XmYB34Z3MsiwJKp7d1PQj7DR8X7xZ40VUdaCjB026Sp0oq25jIJPaeffSr0m8Dc
KYJlfy26rjIJ/jmnfapiYTU0YLPkUu5EtWH4DFFOVJYJD4q34w1htQgIsGFO5hxV
zQ6akzdNJ8WXO+PWaPY0WO22GRx1vHJUWPp2j8q0puAovLLXSq2SOg5++zEjhPt+
XEsstKLa31r/egOmdN0h+JmB38MrCCkZN+v0Unc6inbAggEE542av+rFM7eN5zWR
nhgEiwF2CVa7T90xanqIe0RUtvMuZxv2aBl2D09T9QAHwwrWaw03W7puFeZWKzD0
t26Kqle+vW5VNN9Avgo8EM+H7WJG5/Ka0xNv9gPjlmXBs2kgJsN861KXdGxYtjnV
Arb6G1+uCrte16vhJC4O2s9uvf5B+svdVfE3cDkXNMyyBbcqKCmicPkvJYcn5iEu
KjWFKYVGi7/XVvBalvQW0jrYFe9yo1WPnJrORpKvuBfg7RO6yCs/CSXfkAb6zvCP
YaRboeb16NnQSxCWG3mije4vbu84tGV7lXITpD4yehRpduzgXcYyh7tfpYR+F7O4
0y3D2qI4USszuEYrD8ocg1eqDdcEBNTn2eXrkD+LJUxJoVChpjWnmYZwss5Vo+y1
wlZoGLZnigQHmQzyLOKFqM/lMg83NNqeyHAamhmtcesboMBQRaopj/3+cw2FRz1g
yMeIx3l+tewDF2yRcBkJ43sPdXn1zY8w/IKNQ6bEfrVjz/4bUebImMtpIqCXStDc
EUz/4VFEch8VySsERZtUKuYIhg5KrBn7YOC1ay+Q0dtOJm2/BlkZUB4K3XGDvLm8
o6Tf7Gh+7hnQJeqv94+DtZ/DJspx4TpEv+Qa5JfPUlbaHyTPmIZ4MHKo2ZkofPwi
k2caHQjhnfoIKn96BhWNbTcGGQJiARYs1BFOAg2Yq7cGWdS04tnDIutr0ZUR1oKU
au1NhdX/BHEeqmqvw3dgU7YnXZMHW0ONvur1ZTC6554nH1zMqY/KxZodqFUn6uKm
yScDo89gRLkIwrcbYJHBJFd8HXb8ZNjqNmfeC3RW9vlhvNyVGjdFF5nHqAMjUboS
YuYgLpTlU5NtyiOISMlNvXrNdCT9iYLuN0ketTFZy9/q2QXia6kILS5jugL7oAC4
JKPlkcLpmy9z97jp5ap3InGdOr9s91fAw8xjviAtuaBztTdbk0Q697xiW71KE2lF
GNX9FqMbpM9qln53E5KSVHqw8nIrFB1WfNzNQj7tJ5zK3mkUCUNQiF8AYBYFDnw3
yR/8XgXg4y0zjsve03Y7cMkwGAnEYXCm73eJ2be8jNJdetwQFm7JGqp4fAFn6ZvJ
BOdrcbAi0kMGk52PK/KRIUaBhdcyG0mA/KCV48tHm4cYvFBbYgTbqZNJJY+4Ekiv
R7i5rIepCbZzw3cO3mScvCcSuLbVRkjcJNqc60aly/PxFg8CWL4XUvgdxzp/Zan3
TSyekGVNWFzUAbEUWpy3R5wxIKC/JF18xgWv/Lmr/Gc277258ABfdognIBsYE6Va
AtFVajeWhfMdUQdGnxfmwgSAueSUqLVCkqvzJ/x/2yR1Fa8gpt5yy//mrgAjNJhN
eBURMIQnabEVm8igrYR71myRGibxzebUniYf2Lom/0MzNk4hoB+wAKUk9hWoqq0u
WHY9jAZXjDuDiXXZi6t+HKbXIZJIVFfnLTVAG8NfBlI9Id3id1eimpM6qsdDwsFl
P6mfeW3utBl4huVwTVVXyJ9wi+aBXphGJk5pJQCmAfgtMP1IS9Gb1r/w1FKU3Tm8
WHM+ZNuF5Eu93+7x5fJeXtDoKR2iF+aJoxSzNZeoBWbbdgmX4nYZ43P5ELlbtRcN
Of138tI4Fhre+IgAIiux6ETjKnT5wwt0QA4PJYL/moLO7zpIFKmQrUlHvBFFkkUD
bF2hCKWuDT4TqypwZvYduIHZNijmIX+GlP60fJqmdZoFHktlpN2HgJzeK4n0ZQWX
+gWXEF4QVGcPIY3sveHFb5kTunGLiTr3vySVPyPo1+u57t5R4D0Pb6Uucf8XXGYO
Pu4ZTb+8w40+w++bP91phY7Hf7a1L+7I1jbgnXS+9v7j6fVWBNC/C+BrP+vXPuo+
oQT1BQGRj8MLY2vPoCOfk7AkVKD1qK2oL6hFteFSsC3z11Ax9QRRI1NIiFuBTxCg
epii+h96sIIwod1RVBa0tFLRCf2KN7M2CMVg5VVaw+HNjF+GBeBreJ72xctRw8lN
gS6uQWl9MjA/WW6K0BKBx+pgwJ1rupntElT0Onbw8bTmq8BzCbUtCHGM2nRR2GW7
v+T6cbiz3WfnwpCW3n1jnsro/lhVog524aYntx/heUOfdhEqme085tWN1xWMChGB
N55MDNcFNprku8OcDmrj2FsaZduNATqV6YuccvwN8j3K9Qk+FqEuF6aLKRx2f+wg
kAuFZcvyXIYgLUSg3Z3x11SnXzOyvsZHvKzZBOFBRd3s+m51dQgznhZ0dX06IOOZ
5TRzmWEf9sYJ25kshPfAalHKn/qRUU1LfEqX2hpWBC/lVE1BrRBZRqLGweenXoJZ
g75drhsciHYrxraVjo3i1mzALjqzV9Wq8zJIp7pEcPIUOFekda3Uiy0OmxXrvoNZ
1dUph4UuRY3fvFrfwfyoccmuMiszOdzrWI8z4CJJlLr8KrfOKQKW0YTIdCtODL/3
s1TxT5hf4uAvy1OpY9vtxcEsv93YWOH+FgIBiIuEgfPpcPHo0hPuIzqW6EBZfLQn
u15TfYV6jHqP54+hTZB85x1SKikUq9sxDkJevcbPflh0SeKXbaBjTCc1VWWF/yR/
hVzCU7yYk9ZsOoY1XWdlFS8+Q4O6SgzFXtQyQ8tJszO0b7+PtZUSI7ZEFP6ppfXv
6JIJvw7eIFLztdSj6Cz8NH3+uvsh19ZOrKpINn19afPm10rpqdq+wJcntUt5fLBR
PMjNV2uSt/IPrxZf3jTYytG1g/pmnK+/gc++E9DBLIfxx/5r8E65WZnJatwixrU+
b4fxxYqgdQTJt6uWILjorT4uJobVfq4NV9ON+g4pDXIHu3d5XF2RITxL8UOrUTqX
41mwnteMO1OobXos7gvP4bL+V9bltfp1mjMaBSqal1Acf2mGRq7kP7Z5Zw3I5Fpm
4hjVGQO1lMaDLW/3yFb1um/HQZnB42uYHw+E/zJUnY8B2RhWui40G4K2vA3dkWUI
B7A3ucR8Y493RigfIYJeEyDm/4JyTRbHswQ+DWUi1XT1rsXwO5j4/5LFnwFnz65i
XJaLPLQRF5DVpddUZufPJBqi+WOm7d+o4KadQtCC+XPg6ZUr+GJ4sJeIz7jBQBWF
ttDkVG+l1kEe37k2W8qggCuEzIYOmCJAng+fgxuRCnwcq+x6HEZGm3LEU6cM97+l
yRZ6a5XKTw9tIEebcgMtsdshy++RpsyoA02EdzsoUJ4Q1OeQbvKx04bj9WcrVUo1
qKmUAG9QdpQyHRyOsqwY8yW4e9yvVacjBTWTIDH6txF4Gin74Ccsxx5qg7tJe41X
iUcTiB5Ze6rHBaJEN1eLMbmKSWDcxeXsUpXcXy9Q8egUWf9GEtNZGdpxVtFOwc6Y
5ygd+NwUx2/E54dwL02mn8EAqcoIUbS2OBzeeYVWONyGVWWG/DY2AiCoSzh5t9PH
D+2SqHHCp9HoPp8IAtiCqKzGIWDMY/Xv+UR+gTEtOn1YOjiq3frmrGAez4/kggtd
0Z0DBllgTDbXN7hMRbBstsdU2qAJbZcALziKYN+OQxqVri4PmOo6qs2JAXQVjEBe
NXGdikfx+Qe5WcchALaYpukQ+gIUbkzFRl7Yh4ui9/2WpU5P94+VHq4WK1eTYVEe
1cLQCuU13Pt7r2J9J/Z95lwcJwv1vOmUb8nlZYxu/NIpG1q5DcFz3elmZQxg1FNK
MNfOH3uesSYBCPmlk1k3TsSXCPUHqFStRhQ2B4MOm5A+RaicMZuqttI9b/TaH89A
q1x17O0IsBdRCJMfJ24kGCvFGufxmeVGJ9aYw1wicOlsseRUfOgttoSt5L0OJf0N
Bb9ZrmLL/wKQWm7Q4JFqGAH7V0rhDmZ2v2WRsIw9dgeFprRGHUmTgD9mhmzoGlWr
2WzkW59LtKvCyIA/AAw2wHmxEGWQmQHK5sEuVaVmSMK7kxFVcH1Y2DX+tDCklQRt
AsjLPqOE7Es9ZEPcnIy6XBKVA85Zpd+rC+f7QV6we09rEpntud9J8/xvJumy5dMg
28fjGYGQyrwLINU3S7TS5cpS18uyKncBub+pq0heMmaQE14gsoLpLHEeMMyQs0or
U4ElDEqPC8eip4lIbq9g6bF9M2gpEn5E27lTenug7IS1EDsNuBCRd02DqQBgIJm5
gWnuRAuQIwT0Z7+KsB7OhnVVNqsJbivMaFVpXkiMgJ1nNDB4dbhkK0YXOFULWNvO
Jzom6yEb3dztH0oNaoVJtHJhrk8EHvd0SPrNlIz+SVxXha1qO228g/mTL3+it/CA
dYXcYx3a72+oNpotlAv3pXaIaicM6BNMkR2dAIQVh/ZrTO3BF2Irw3q3UEX3scM2
QNreZQV35yuB1RmCCquhn4WlV5o48aC7aW7ryWjMZ5t9Agrc/uQdCrT+CofNscJc
o2TQZ4dc/S4BwgSI8nCS0MFbB63YNslEk/uY1xYoUYL7DrgWWbCzyx2EB+HRocoQ
wQDBcGa++jMz8ivapC75esUIzGH5aG70/bnHED415Z6fGlOqZTRskHH98fhRw/FG
Y47cnj8BLIu/s78VaoYbQbpZF698NS8/t0HwGp9RZ+c910XBn1bmUf087urn69lO
K6xd5IhI8iXZdGQ0siaw4ppjLmJdNUAIehEWpazs0S7Y/dFshikKlgM5UGgGTm73
LsMM05x1+FqZJe4OoJK1+L9uI17DQ+mrYq6RQMSNM8blnK9xVOU9z0/qq2z3jVrH
6ekXpDBY+l579LCsCc1oaxD+mnFqOpf8kd559TLk3xD6eHrQ4HHCbVR43BMq5SR4
Aeu7pujuuovweDMQ0XZXLSHY19Bj/jOGIJVvH3u5GiJ2PNzplyjP62QmIVodUl+9
OQBNS7YP7M+8Bw85X51EJSWJSL3ClqSb9FYy+CEQDnki/+ksIvyXZANAWBf4/x+C
DXDcR0qwQOYAdaRxBRQutGN+2jKpK0tGcqAZyMbzXDpWEAcF1FOyW03rGLyNdjf9
fR6vqQUIBhiDeP9nOrx3sXsb4dT+RN1smeimPSGEF0BfSliYKOkCXV2Goh6HA44S
RbDI1PQTz4gPYhgTKb52o4ivZ06ziUtjzI8gY82YGMtBG1CrSg+yxfThI31jNdt/
dD4f5MVeRzEkr4uLGYgvIyyf80IIPz9Al+qaXGzac+iaKoYGzE6DNcjyJzt5EKSt
e4SPIAM4X/X6ud0DiSuxveFbtqW5IRDiJBq7YeRqfUXbgqkJUhzuqGn4aOPjnQ5Q
m/feJVXOxp2MIM83L2liVUH88WYwayA/3GTH4SxDuxZIFAlAW/gddPSqzLxWkTvW
0CZEgKc34i2/V7XFl3LmvsSBlADDmeFR5CMwNsOqT2vV+FGM7ifNh6HmPtfJ03ez
5XcIiIpIdyuBehReunAfHLqNO/Ikpqnl5duTWU9uoYThHI4AaycG9kRkRsqH7hcv
NN12cMbdDMFwee2xu7luXjYc8c4hTJJmp87dfYpGXqhoRRkLY23cL2av0/Rgahet
b7GA7bkRYC148gJGFHIxT5fMOVw9FbAEo7YbPfofrZVS7Hh069gSfn13K8phNA3R
nwPVUCa/GF/6OR0d1otivDniQkcl756AR96fdx9nqLjtY6zJCiTA1X5gW0lC3Dj8
W/PlKzysSj6BFKe4GtcM6yZb+uHjk/nxyccR7SCmfPf1tINudcldNK3GnHhBPnOp
hSTitV/YlzDL1noV9drFE+eCjTxcrVr4YklGBF04RMIeGb840CWaDWAJy9IIGyAm
5DbJrEI80fQ19KU/GFZpkqpqo63NxT0bzV8FfDml+iAeOQPTS7YN3LjeNadBurUX
FQqxWreuPKkQRwDp0YYmtar7qR/A+v+MWX3hPK2vXlDT/tOhjLfZ8vZxtyKGEJnz
EexiRya6gQ1uO0cbifvjpjKuo6bHlp1KZ8UiK53lepsB1QjXQ7EKBqef7iSCAW3A
LsUepUZxNRgW+ysAJ9KuuXGjT49eyRrK/OfRHBG0KlDKj5Hb+ZpW/Jo9M1YB0YkY
1d9oP3bGG2IF4pv/7/3ReCWc6F6dqAst5DKuel79LujFdfLS6jZH20KAbl5tzcQD
6TqCTsoEsdxAq0QzFnydWeqTEvU1wAw20QdU2zpVnZ9ICWunbuu4GBKmrWdJi6XM
AXniTMoI+wUxhlwcXh/88I66vDkleYQ3HDlYI3pvP+U95FEl0EKIpO2Xm8A2YM+J
XVhqCN/jo1ukKIMFRzinbn9hn0xR0gq2Z8Ejn3rJQQQaYBEelxR0qDifKGYZVzx6
tGx8uEu7OlEIgKHdF2Umt96mhjM7bnsJbGKfY+HhWPSfxYKE2dLn3+Iqq7yAEPJw
ym5W3XRGaUU1ixOIfrE184mYfmT4RqV497qkNUlc3RJ/59bNIbpC34ZgVynnKxjO
5+f9n2g2aSdr5XJb7PBQK54+1uU5N4h2pvmPLIJc3rP+XtwSn4NA5SMEZeCOdyWU
7lRstoyW6Il/IceB76rb2Pg94L9YRDAX9pux54fQPsui508ybxrf3FruwjKcdgcM
9PAM6RryoiZxcVOCisd6EH5ZL1NgI4g7Vawxl6oNSWjyO/olQWVrij4flUUvT82L
hajbBchUVwn5EHkOidgW/of8rArRe2XRCDP0YLnMWGGZGnA6nosrYHUo8jTdJu7H
pLaLEKsN+28BEejYFuyuEzF47uRBuuj9cL6kbX1P8NBaD6hyAGQyE1P0LHH8dxB1
MHkSbwMKZAIVWF92g6ZtJhPzcaVgh8UYVR7NhJAD5FKQR4pezxHqbtCE9DqQMGFH
oTYQYTHRV/OEbNP0QedUkuPwP+8VKntiBY06h9T9CBffzRb/HXzGOOInT/UYYLDR
78lbd7kfHyBL+XrLuEBoSHH8lq0V9EMBtbU5E1yMEb47fEni5Ojf4UXIbAxU7zzs
KDTCPtaZQP6WN3OwKqNaJytTzdNw0Kze1gcSsZNj+zXMrb8ML7siZLbSkcRxEpi8
0PbmsU0EgZuDDjC5iCLVRMKz3lCLnjEM/XEotDf2VWbJbOg7dXsjiazmAej2aosV
TDvdEHmEgDZoHwzc05qoD3gIUIhdJJUBlsh+zAxqZjPcVYoKsYJK39NXgqbCpdHU
F79ktTS/kfaRXXTBmEjdKF9tAHXlPGb6HBcWr3bcIJtUXTSX6BvrT5vBJV8p5Dq1
eYq/smgyzTDskYqpruVQFhRB3q4eBjkZJpYLXMJk6WsS/0z//Y+zmdudJeffRw6K
Fe6W+1mb6hW3vK2Ew4qkHtLeWdu3ciLYuOXYKTZFDjUxtJaAvXghFPBqbw2Y5cjW
XSYUv1mVBwVzEs3misF0nZNwjZ1A3WriEVvEzTxvOsdAULr4NniC1YrTQGEd65nn
xZru9+LhM3uFokxO92zvnmJWPC5qf0XWIVnjRN/zNv0Dk5ZvQ1uEOECEA/wQMRVi
pt2pDovd9p5do0PJSGO0TDwE4GWgQDjWxL6dASvQ4RcBBm/RGLUb+TMnIgLbK+1h
w6Ir1lkzwm8jGbph5Zo8E3IUFtycrTrmeAgOEfeVu46gcqGlgRbCGGd9JpSCBcYe
PY4R5xffF8jEmqQhdON+ACNh3XbkBIjBfEn11rJtXDFGLBmogbLpMKKw8nWDfkvf
J6eQv0pD6sziTD7y2EWk+9uZitUATDgJnY9n76ial6NfS9fA4NuKwcBRNtoE+4gG
4hqHpy2qwf39grJOgpSyN+99Fju9dM3RAEAThB+GyxPgcyT4WuQHRfz0KkUnEDfe
WcJHuVnI4WW851MOOkulYSOZDvd2eCbchW1+wx4ESeYfyci6SVLALMQwm3Xdt59/
LeZPK7RuAijhsIK7BUDsrwvGTDB2h4+5HbDxAzLJ9ZXkE+eXJZRfwPYmbOKc9Xfg
b+lFbpPjSY9olS7863yPLuiCo9Mo1TFScifq9AMUtJ9Cqxng5tPXQfq9n0IayXtq
57yQqk2Io+Gf9zaeKFC5DFqha3A1iI6sJcOseplAe2shlaZ/5v9SFSf/nV8wsFAW
qqGEUrduD1fcvd4cU2964vKOlALhufWN5rhBTPE6uTOQzY13AmgBFITBW1P1BB05
j3pQLVQgv6g1PA+qZdG5HKHpWU1GttNpiL3aK2HNpuMli2TzviGjXErdbEkaK+6u
sj9jhmPvlfVe9qCBCoMlL16RL7c+gaIV77vqGHRwck/BUvxUyKREnE5QHovj1DXO
rhBGkRaRCWW8+ENXxsatYIn9TFlYkC13EdsaFbi97rCCuj7k/aFlXQRqgOrCdPRv
9qy2ZefDLuRvbgm17+nAdbWezQBYc1l6AMBLQ8A+VAfyZKVXn2gWV/8XLCUlGP67
YWu6RXXujvO408LqkjnFze1oYy0ZECJxHk30ekmj28Y8XB3Bj1pbLOn/W5Se52hf
QG30S3LIju0jfEjEZfP+nXBHDbzEB7FIV3eq3y9sA/badpLpmMOwB14mOJDc3G+h
xbuvAXlzuJ1B69/0lsXsASASWAdoMsrHTEFOYz5ezs66EWXWG56OD0ot4zZtXqUA
IRGK45GPF3PNzsSJQy2xowIsqNBdzQcnysKnIPPDW2CSKQOVSbGYMFH2Lq1YxT/N
Y5+BJHhQrGPjgM9+PVxkDdCdKGTde3DiV8ReQ2uxiHBtocTidRM4ycGIp1Dxvahx
5mZpBYHPn/t9S7m9W5yQyEkewIyFD25IEJnmJ0sotbt1sz70xYOqjKtlzEVGe9X1
Z9Logmisw8HOikth1k8wu9KC3oGMPLg2Xe+a/gXKinh7JA+zE65DUQIhDt4k57Nu
fHNgxTVXhs5eh5pKmBcXdsfEB5QGV6RZrxHbx0uPiRO4wh11H610YCJhJiZn3teE
fzxS62Z4MsEYLuraaJBAkUGUiYQ7EMsoo/qJ7lZ3w+uqCX7/ISFUbX3i3aqviAKW
+GzJ47T/nz6kDR8/+NzrcHptCS9c6HL7p/2g7SrrAlTGy424xzjbrtlBhLLr1/uI
sdpsRFa7E374noR0bAr4gRgNeJj8vd+FowAx9oNcHWUS/YgflusF+4bxrUJBE/eW
jywn/P/9zTerffKjXcXWLFmC0Cg+6FeRA2HaFYR7rsiywEvEtDOClApiuxdQkIMu
5DaORWBWK0zgg5mFGFyRsvMUoZ/ziO/IW5ZhqpJy+ybwwanSxu2qBMj1f4orJL16
AHQgDaB+eXstP18yn2Z9gD8GBXt7BWLqoedJDf550ZledxBkXE0XwI4FPQ9sdHm4
szs6joVer9sJAzzaIyPAiBUEtbCVAXtGE+gJsHhYHTvKO5MUZLcXYIFbjw+uvXjt
TaxJUBzBNsXxekcd5K2hz8D9Rf/7gMGqpmWrTtpQNzCoQGuODZtNM5BRQkGXv1el
faheiO+Qd/JneEEGWNsA04M/LHJFwNPcwGNiTKLw2yV0En9lHwyAwCKLs9Dz8O9V
by1kAZzI2caaQipiZR9ATV5jndzPa2r35tfHYRNoDgjQTr96jAAv6vdao8wZBCDs
d/Awd/nVHEeJTLSO84sGz1h01ZnHFauyLuf37zVdq7WsbJnlLq+oIWoPKenF1DSg
is5/p2JTm8TABWl3NQt1ou+Tm1qAE04ZkWlUmPp4NFAKpvmGwgi3YMn2+IZvJiPr
RxzWMnDYNfeSjZKUPGsBkrjFc6766a5jGp+kVTqE6D9artgyyYoOHRZ1NPTChveC
/+JwpBGDWRjdZ/OuEQAtqQtFoKtA1+SpTJ0Aw0FSx/TyYKUQH/HwTa8pv633QTEX
Fe0brWKvMfd10fOig9tK+RTjNklJDOMJJ81O0Lg7MjfeTipoZDpGe1M5l8DTT1fS
3ilaJ1wO05tpWs+iabENa8d+bXN6DBD5e95/u7Dq2diBl8B2WK7v8xY8Vl7jhS8S
mkKEeryU60dPn8iqH+ulKnsJtzs/6UDEtfyThbSo0CRzwybZ4gSuwaW72SD5OLGd
86YDwlWTcygQZfBbdDPQ5B9D2ozkvQlWw4Q/+Q+gaL8yqBDbohU+wsn5u06M7kmX
TrkCHJxr9xTYTtlahW7Anr2JbvsrrE9Wpo+sOTRmEEIJyL9YWtIaxAHs9whWpBMF
+hgJQ8REYJK/Eu2vMLKulZBoxn2HqLUJ77pIcKEdMuHOQVcrkive84Er2Us7dw6e
3nt2WNQqIjjQbQP2DSCnEL2RmOskCxJPTEufBug5T2cXt8mibfYkGkPR4pOyl5Li
FEQLFl+RxjBc/2RSbCmvqYOxP/oV7L9CXkf3MYJx2nuGwQ+1TpnsII9fCOX1IGIr
/DBCEaPpVBw1At6YtoE/Mu5pJO+s39z7srj3mbycoXFYjGBUj5sgkI/uMdeGAXcK
7d0DnvyGDgfniNw0etmk4KrG/fOaFzas5EA7w5JgaqSVF35bd9B19/14uAnwrYtJ
q/xil9AwPaCq2jkW2RKWpFXYgJBl9WCGvenrov99MHdltjHiJsRJh3zYuvrmObgP
RoQlwtNzFoogIChF8biIK/UO3qtmWIWpk1dPBkyfEdPfwe7INPwwaMaJNHMfV3xd
0r4VrWMFYaU27w4L6jf5/xlYJ0yNwfvvYklujgdrRCiQIcP19rsBKi1yB6ssk5B5
wLaUQFvG2qERvQLjpSPfg2xi/KcD0k9nA762sZPg9QZ72mUmASpBIbvCxtKrG9yW
qwbbSVjXB7z2IwTL+1v51UO6Sb8gCK05Bjvk00C6Mj/C04KelHBCq4KGoiVFNYof
XNysO3m2WwadC7Ba3V33MLMrlI1ONi9iSf9O39VDak1ytLhCqODZImj+A/fYg0Zj
B39IAxVrrSzZpwdcDK2SubQMohMyGvb6zIrugCfZCI7VZvwINnIegETZTq6Ccpmz
vMn0fxBQdUh+mtgK7i/LXOc0aii9gcc5O4B/zDE/3qhrMLONGz7pte9ptZ4QgG7l
4UdcTicDR/fgq7mskNmI5SmesAem6W3ICbDD8TTeXmfN21oWcOMRWY4YEM+H3of0
I2E3cZ+rFjbiPR+M6m3/O1S2aLrQYn1rYCiiLBK/ybWX5xuxilYecHpykcadILZp
SiAqC5sGgUwUSFtmvyHfuXpi+BwH8tgj6XVonCFC1fXe4GR4H85Irq2iwFOxY2hq
TW0ybCsMUTfcMLzfXWAg0zCJP+4n6GwFeBvuGvoumveE3qCdW66AaKAPRfoFUgSN
Xjg5Eh7ZtmqFgfML2RX1NZRbSxi49BYIJz2eljmitSVf29eVeMZezBTcLCa55Tm5
dJiz0Eh3fjip07BTRoR/zn/xCkzW0bGGraPL650pnEkPoLAISd09tlossec/XK6w
GAmsPHeJuOwqmwsYAUvg6zBfd+oh7ZYsrzHd07wrclD0wN1fDIbOIwoxc3Ko6ItN
WxEfTC3N/RLivfl7WiatNpGyzWRj2J3T16DpJ1Eucx/Za6+4hqMs7wT6RTTDo5S5
8L6ySqMBRUF8KlgSYU7yUSHZZ0wnbeYOUH/X0M7i7H3oRWCp1JY6OdRWZqpWJisG
ogIr16INW231fYijp4uqJkCHPXapnlXVqN5cKnHOqt01W104nuA/T6jNmWztPVgj
CX5Oi6TeqQ+uNeZOsWwnQKbj6ZpYnF1ALLvV1gvqVUh2hUs42OchCAEJ+G+j7yxl
GVA4Zkc3Fj3Ur3k6a7gyKbeol9f60SNSWcfTAwUj8ZXeQ1DRrYa/QGyuOH5lU7YU
J7V525NUyn/zQQAqJLLFUEzfEX5Xa8S4gEy8ztvucJpATLdGRN61Ka78MoG2mnQh
hwr1LnGwiqN46SoKoWeTgHecrmQYmMJ9qLJmN2uhwZWpchwNl7D9XTpO5c+fGrfv
7qXuZ1W57lLLKMYSO9SAdEqo8R4YhDi8fweEGkTV4+zqNNjyf7EvPeupbMYfC5Hb
CtdBE2lQ7bq9JQ1Iny5ZMxBAnGxvZjcd1OkSDUF4kBuhI7hkEKKQ/c2ZYtjSw08g
FqWuBe4vRkV5gIyFqWfRwKShp5ElmAFM6YZkeXp+3mjecOuZkFdqpPjzAheugSik
4C605kESLFxw7Ax9jfBpxHihXP/R9CMBx1LAIFWQGpdOYkWQfQKXgAmpF3rptDYR
H5hhBX27h8cJAjYbXBg1ErHRmOLR4i+AWwzf5Ut98WbUIacOrWMi4aEBBMDIOiI+
moA8EZOzj33tgqSLOVI5tdC8H7lxGh2KmCWZmLxyF2VA3KSdkjW/+hKebMScqdT1
bwVBMATXLg6K9TkDXv05vHX+9udLwDRSj3YJ43uIuQdPXmCBne3DuvkzU0UI6xiS
hmmOYdu7TDjdwvSkzINcOcuIHtrUCSb572HH658hVXGBHksaqICCYFPoZ52BqYuU
UJJSTo8b21WXknFPDS4cOTnX4f20wsXbz+7ayAcSAIR7/e0buwISZU0tVNLCKA0s
A3lz0ZRT6Xas6/rfO2SrW2HSfTzRkpItcdjOAOIQW1Q7+UsdKDQqzUAwMbwTnfog
7hajOtiJ/h/Li6per6QGzNBwqUlLxhgrqSbrYUFiJzzYGMawJC6DFGIMTzd0mDCD
e7iXl+Um92UbmsgDGtKobq72ojRe6ybrkjheZwQUVXY92aiA6hIOvN6d+Hs1g8zA
Vh8QRu60faFKuiEdQkgySloB7Ng8U3ggCMMwclXcI8MsgzVX+xShhN9jOMNO4iNz
NdpzDe7zSSBkt8i/RGwYmCZJRzywO4RRPdl+Wmk+b8XNCNUUD7hRNR2xPHAjHTWG
l5V3dngskULCFctlaSVQl+at6oG4yaGTXzj6p7CVAYDVMK4YbP/bWvpgNnUQqC2i
ZJ+4eP670dABhxCf72npOKH5twvdhfEqO02WE5lO2J5vRKUTfVQtq3IQ8CzDAEox
+NVbvZLdYD+RnNHhu7VySC23NhKpZWXVDrUFaJm8EcLi5F7Jc5pbNSWcMHJr0QAT
i0wO8uFcdntFf8kMa3VIWPCSaIrHoS3GkoDHC4FMKDtKNKuIu3w7Ry0ouhpiTK4p
iLAL0AUhe2cZnIWXjcmAb/l38j7p+STvqHHKghcZZZgd8EQge4W4J7+XkGMcLUQx
H6Bhb6DjQsnQNWxO09B3P6rSZ/V+cjLCAPdwUnmfNoHsRU/o+2HFuJvbhevVTwwG
0KWttuTBTNcEB78z4Y7mrOb4TRe/wtyAyuWDtD/gQPi9IPUUI3hpUE27P/d4jpmF
Pzo+qySbtufKxtfjgwTN4PocZrbXyM/y0t5o0DlS++GhgTi+LJW0iz8ku4CWtVdN
xClXs9+XjVqBeYwd7RJgMCynNV7OXfXWb8RtmUA3+v4Or1+FcvcQI80qLqkCqeqa
YVkqipmR0aMsWl0CkDaM5UJp/jG1W0oBvEpsKRNmwDFERELa82SaQe90rg/9Du4N
LCSY8bSPtW4EF1LKf+qQ6Bs//rj7cgIVCRG2xgSOP9MvYhFkRw25ouZA6hGbAjA6
KJ3PjqWsigpckSSkGIttDO0ZYJOkH1XT4jVn4TFA1hcqjIDL12AWEQu2JNQHVKS2
dqxGnRjruzlR/jLYwhJQlaNyL/AmcbfzCqckEM3z1xU0uq9TyR50++1PHCWpgU2g
eOCinGisMHCbGMHFP3OLMFzyVWo0V2VjxwbZWKa6B2IjSva2L+8XLTLorvrSnSMs
YPNw8PS3mM7niVDZaRFO5i9b0qD5DRJrj9Cn5leC/UF1ymBaQiNqOpPHruZPpl0+
JNpSdmGMhh34nDhq/qk4R0H/vk0AJx7D53jGW4pSGKoqh5mWQXNY1alacysduo36
PxUSdpfXIreW4GZ7h+BhbohutnyjQcKtS43ungS9VB64pLL+Gm7fgJTynnE6yjeu
jPWirBdTvWxFYEnRwC+a+6s7SHh2IqDtE1V/1vnA/4GKle9TbTULSTq+N0bGddF3
8tcED8TiguAX+McA0KGF+4SwxNDbfLE8fsMoG4g8aDldipSx6PkB/3UUqsIVXUWY
cRZzrjXgFW+ntuCW5jrnZYs7BxbSX35C+HRWaR3kxkUpbjUByaamvvyUXg8Y8RyS
qCpxuJCidSDELMUIGGH5WBxK5SXMCdrkcV2oG6Oje4C2XtxgYyylgaEdj/T/XyXx
4ngP/J7gm9THn8P9oY5x9/lqJYLN6+5zNGkPcrZeK0gA50FOw6le382yf7+hgov8
008pJKgM/dXu6T2NyTB92e2bsYc1VHuGAR8jmx2DeNFVd59Q9oIzpK7fj0/Gp1t0
L3BVMPiNgY6XgxWMxx7SVMiuMplcIpUH5OSx9yuCsSsvPotlSXw8EZxtnb3kJM7R
/BaYajI+wjFb/23HqsYfs/BgFw1wmy6zX8D/ixMW7DzrdbJfEJ2abl4sJtAJFK26
5qYFeDLQwfphqBrnXCMVkRHwHPMMZ1AT28NrgkrpSii9T2vehmxNZfB6UVD82aXF
e4LvrI20IvVR/h7gptZ37tdQIDN/FaIChY8VBo90kOBM2oEJDBDLBUBjz+MtH5ap
TU0yTyNX8fQJyh1JkfT1FKBal/ahk81qqxiF1JVUdf3OZ/3iiht8ZMzOPhRsOq0+
hLkTrh3vCALZ4vg76Ku9FEAEo4ZuQAPgdl8eNZFEqXZo5tXi5J6JwuHxgYrupMeJ
5G2/cqQV6d+BH9i8nlI6HNrnX5bFWhBzm4RK/HB+lTYTNGKQpeYiHTiQWz0ggkFO
u1r66IKPlGBX7KHq0dWLYwi8Ytkpk69HRcmsECppuSsh1FwTZkICLbd1jdN79hvE
jpKXzkLssAoAbazN7pq0a6jR27EPcSjz5v8Ry3ZiSgfG4mPj3LZSB84nBOLNS3PM
c48eTnipqLbbbkj7LNgpXYRqbtl267yWgjrtZHa1OnagBfgIhuY3jSazDuF9idh/
RPqSQVOysxmDUM4Qw8vd7tB9BKCX/ftZ5Rg2FDn439c9YWMMeWT2BUlJ59wfGPcu
2tB/W0m9f/Kqs1i2p9+GukzVNMFgonxfNmdfWY4/Ang9/wS2SW2T1mQM1AKY14cI
8BL9A/ICIfEo5cZpPUlwI58/qZJyR5ZfJZMp15aEkcgGWY9XRQ0T8Dx+oLzf6qp7
FQj8dYeC5IaJgHEEywvCKRavbiioPdO0mR/nYI3LlN+MiePunCl0Q/4ewqltGrkY
6DY3eLUeoTajzbvBvug2NiGS9CaW6JZbeCzY8o5dCK1V5QbI/omKA5VZVOv+uNaB
4FsdhPuqI4185XvPL/FbBb+QOmw8b28n1e1QE6VmN6GL2FW4frDnDco0pIRGd4GV
Gxs+LDLMWFGT72gAauX+6wSrEvA1bHRUV/C2NLs5nTOZcO+nHq6jFErtAkZLZw+n
xRDl7l+Md9bAo/2qfxBicHe5U16tcljn3g2YPUr9nATsnPaunvze6J80EGFUKc9/
8pBCsLyztOKCYqj2zTMA83lKeZcruQVAmqwCVRCe4sMsJp5hCkv25wxY0f9VoobX
1AyD30FA6sdyHoNliB49tGexfR4g102G6dXkrtzzlitXpk6oy98eosn06urGJWVe
DWiyukscH3glH6Dwgy3varG5Le4eoZsVu5obHiMGd6x9uGpGHJRsKc3E1ItXXS0y
zbshhf7XXVD9vkdLd8TJcVqmvMDCTqYmSuiNBx9c/E9iyxFADp9wHhZs2weeCz3f
yIMofuBFZq0vE/LCkIsKGrejYIKSCsEBE6KAdDauVmN6ZgB1Fw7j0/9+pbxCRgxD
qU/nOkOCJPbNlFf5cXpJwwkDRyMlZvcpHm6feDaHrxV1A0Jjx2EeeiaZr7X3epZv
e1d/X0GrW1mUKrvIBjwKlIY0MpJyNw4RzLPn6MFRx4On2qUyP22QLONj8urJTUz3
sKHwxNkTchy0wJwBt8GcUjAveoRaqeUTRou1UDmteD7OfcZwpHriqcw7UE6NdtbS
gZ1PWzne9xCfeYkEwTMxfhKmAVQ1tXke0ffl/UW1tD9bhavubUreIzu7JlzFmWkb
ceLpw57W9Fu2ivFth5Nzg2F6Xn2BUt2FoMVHHGCaEMAHUc4yXIZdJEtyZ+0RplTs
aVGluBd5FkL2c+FDdPHz+b8pqzoOM72sKLBHrQwLmEUcicf6GqFGjvc8/+EkubCm
BrH1EPuTRRz1uRFti7YiqPDTQR7UgxAlfF+5/7HYL7oNYLqkfW8YFZYhiT9dlqic
v+oHHG08aI8AtleSY2DKGcT+FVDLGrxqt8cQh3Kn/B3xdih836pTFTf0fWFI+Lna
+XZ4GRFlD2Cwj24VGC5aKvtH9CqV0tlQ+lj/iFgPRykN1nFfDzqENYa/M+V2WGwi
IT7Pd0nZs7IksKWc2e4MRnqkEqMQu+49aco1XIU6PgkyR+cbPl3C/2A1VLptYSpb
NSZxs/C4FbhLRoAq4SI0Gz1PLWi0iKwwM4ZvxDBLivY7B3Z+bBwu9UpG4AdyPYqs
VFgVAdz/DXVg+J9TiEkk3leEanx6SJIHRNuQ6VU/tIEOk5/ADmubg4kpPYaIpEiF
1W9S7pvSu6VJW+IAaZxs0kO58ZLjh5oXo+HffD2w18GBNByzWSi7ASQBw0lFQOHt
0WmCi9Kv/FGGZqQ7DWtmIEiXf+frtdQO8h9lzKA+O20lEvlVaj3k2JCktxXgan3U
wJymzUf4ytz8udZmcFSRJjmw4LGqJBCrUspPVTAQkfWqRMH7+jcNH7+eh2C2nxky
mxr/3jgKueDW39HlxOr+cbaIw7QWm9LbfchKWMk6KNIK+LFkbu58xc2WFyeOXq8u
h1jI4kDxbNJINkPbUyINNiC77MVua4PA6Lks/D8K9m+TdiBISLbSlS7V97zw4S20
it+yQPJ2B6QFe9NMQp8V4kbZyPQP5nMubDJ5eDsRsZZArTusUwl6Z4oM5i/1Fb79
3twfFX8bhdC+f5bTlx4UKSkunrCAveGRBKQJhpyDUDAgNXP546VKkM/TWCNAQWS/
wHLpQSSUNWzfTCyksXLiSviMmckJaC14sCrNiIuidVmNBT7y+ly6ta/nuIHWBR+o
2+f8fXh4B4f1DmpwO84CbMfWY9XmvS9MHhgljdExXqXs0FzYMck+a/g/vaOOBvU5
002KrW2xowAFPwT4kBSuNwxaZK5OhljMCAEWJlx4LwfS2Xclnuc4/sve2IPRlfdH
hXwZq51Mo30DwnCZG/+OpFgXTYaEM320aReoJN9/Y3ipw9LVXXB4U+OXLNAb4k7t
iv67lZw8menl8qSe3caDE4KvnUq7y71s/zQ6mFYEyPMhl2ozWfrVdFcmnPNdltQD
O59Ix//tbCdNBV8/KviBIoGQpFkjfzdqH7182IUy3F6RbvfqahLyvGyCz+E5Gud0
po35oXBGeF6FLvTMz6IliFKIt9H554S1tnIxkb5ii+cLdRgbdL8WIdJQLSqQfMWm
wDUeISeCvkIktOxcDgKFzNJ+CpJ/AUU+YJdyyY7SXDHv0ohTgANaaBui+Umr1TtE
fbcVDXBKcSc15CRLCg51bzuP3rSZvG1rIqOirKxrLvgA39qlnBp6TXYAXa7iK3I1
uxaF8JevpkuXXYrDt1DRTgWPXCAQbPZFSZ3Ly5QcU0EIv08JBxZYCdhArLGovhZJ
LjA1bTwAz99aiX1zRXmSc+cUL9jkkyZMe2EoMC2LA4mNGG2IclOEz2BxwlZ7d3lT
k7Tc58VQ+2QSvIiNwFSaY14Tzb4XiotT6JFYHZldnEpObnql9yaHH1qjD95ulTPp
rWJVQAxT+KiKSRz1Y0DNEHfBgDD8cWVghIiG1cB5cQmyzTiiD/ovCPpQMZDFYMVy
uTuMs5gGm2+aqugYTbZr5iqDyz9oNo8framxx3uEDqSeGig6nWcXtlgkBiSydBq5
E0CFedQrXQKlrft13uKac2RLQeepG7/D7avqQFIiXcbPlvtj44TfnqNrXSx+N0L6
t5GAFVQqLhwmXjOsHDUdQaTh+IYfH4Z1k6V3G8hrKh4QKPEj9/cub4R37pQs4SOq
qwPtCg6Jm7XZ60Lu8DMH1wxUK+h/+BuJya2RBdBVCQeudniZZLK4bgqUoEpn/9PM
uOpvJKgwLiVUtGLa/ZU3v9EQWFcvchcMpJqAu77xMDgGLxjtDlMoNlBgiE+iisL9
mivvCdUIQ6wDDH/ZKA5khwulxmjfqPefCZKmacXMKvGXuliB41wE1K+BfshFiRbt
qrERFmD7G3XpLbFTd1Yup4kUcYxRGz7girNTnJZoiVNnmcDHRQe4hKyCmb0/ZIaH
Wf4STXj9ORfqKteowyWMzJnKQlK7wvsJ3llBhlNYJlUF/mRE8K4jfYbtOMPn5SAM
ZxpF1ydYrJ9P/rme1xvAD3aX1fCX79O2cZZy1WjoLr1QPzW0TS8SCAYbWHKIfvwb
zkz1BrcXCZihMI8ltUaiLnyTM4Xfwm6l4/3Sw12EiCn8vo+05T030Du8wrhhLdi+
J8sLFD2KHo63iH0SnMfkL9wQh9js0w0CLCDvo45R2SBmVb1li5r7gwkvQC/FcF0g
OpcKx1YYoGgnnErMV6YjS3N7u84KfFvWmXrgyK4j8Vf8pxildCm/1sH8Btb5huis
LAjljZveCtqI8pUQipP61aHzULW69TDm6C4dT0ZnNNTirFuivqkA78MbDk9iNgOx
YrdC/2I41J5S4KpgucTBUilsVWFyLC2s8OXVWe7ZMZk56DHE8Y0llVfqluBn6ZkF
4sR1uQzMU9IstMf6ruEsguTQx8WtHvYnMi1jNDyilLoRjrpE7kaZM0nq24lQ9l2s
1k8cybufq+TwO5DCeHe3oVHH/C5+WV57oAnkOvvIsfrEX1xBwydjHRc0tKjJnSc3
8o/R3ThOHtQ8CF8u6Y1aR8SKo6H5k83NmPa7KXyqcEuoCGSWt20qUorMu7FBDENb
LDdk5aAPASFIklxqX0ZDpKXwxavWlNE5GjoBicUQnjhAQKVP7jWVcdSQ2fzuq3/i
xcmCgI/t/D3OyJfuthk1HaeLZCav3642tsb21fJq644O7Pd+vOeDgqJGU+5+hqKU
QUT2QSnxjCXNee6/S1tHafbr87HY5eEkXWDFYbocb61V5E615hF6qGcAuRQer1Qr
F/WCAKlKkT2Xta+oDrjvj/0vtWkLtfxjm5S97RBMUYNCNx6/mei9af5kNaLjthzn
TJVDpX4TUw5xrZDkmFJiZt1bdo7hpb/zzkPhlhzusBjdX5euG51IX2Xupm4WlX/v
C4RFo7n0mkcNpWhy2ei/8hNQ1qDLwWMqLTzfMoDRjPkLFDiZeFw2BUv1vQxp1AxK
Y3exFzS219CtfDs2kdR0W9y+jkuc5jJFkgzMBGqAYVrGqexSPXhrn0vTJT6ouTjy
yNTW9IQ954efzSTd4G/2xjKn24AIVTlRHBoRamp59ODyxzpT8va8FcrXwhj4OM8V
x+W5jF3/C+3rONyFPlB0JK4bXdR9rNCwibn6rq4mwMeuOG9VSlPdW1+eq9rgvClV
UtgqPalCSW9gLE+CIbd69ZeEmjcsrje82apLHqtjk0zv4BIwBWOu0nWmZctp+LH2
3SrpPsXTHOfQOB1Xx8ImodptjqGNocz+JkTCQsTUZ84QQI0HxQwz+6H3UKUDMRKq
ze3h2UKwGNPWTs07B02VL5edFReFnyDIlcWIThkOYV7QS+kFqraE1zcbDF5Bdb/a
XY+hZ4r0QUBH92oL6zK3zoQhh4QOD2+XWf85vJM55UXYj+3sJ5/sK/XQziibRgaG
C+vwqF6AYkZ8+DsTudPmDpHMDLcpsvDOGuMfkS9PzKvT7x3f1qYngJAc/iO6jTR0
K/IZm6Apf71px0uxY7c9hbB0D0UmM8PxMzuXdqv1ICds7qTtglAkvlVVakJEBct1
EPMoDK0mfpBWvRo2sNCkdw94MVdIa1zot6LAumRAviSNWbyotlVxQuVPu9NT6B2H
lPNJT6ljEhhz4zOg+b8/qLlP3pa5f3VeFY87AabScOfetepsNcatjFVTo1Zb3Xco
mQxIFj9R0pNU1QOAUwnbe0BiNGYhBrQcN41/giOfc767KIxiiNrewwGpR/7OEHol
XCePoyrGzXEog9/lxl5bATwz4QDwJKFbBG7D4Phd+7aOA8jLhhGriINXr7+WviWL
aMYOhj9MF7TsNllV7oqWW7LwWhvDq1FBXT1zGkK7TYlE+ZPslY7nOw0+Q2OvqXgD
yodM5YRP9y/QT2Y5AC+i2qSt+5r75uCy7uFn9iqVN/+Z+V23yPrlnr/C6jqrREsn
YsTELNir5NlqysLeYXzFBap0vOZ6Cw5rdF0NYvGwBPBphdYQWQzmvX7cRI9YQVK4
ef1/UbfM3C0SxUk2rDdtK1hv0NG6LeISVjQvdf1pbSI2DWoicxbQsfu7Du8lpUBA
IHI6rq7fYkEqdP6dXX7qAvyhJJ6gUwxfIamcGroNaO95xzQKHZqhNba0HTL9mZxE
zp1oMCAK7dlsX9kW7Bg8zFAi3Su9zF0bxbDL/Nv6H5fkiN8O5HD/+tOEcm068XSh
k2KEwnqKMzGKcgA7MD2NVhwGzr5BebIB+9tUPa3oHLhlApSOP6mVvvXZowWpXvah
yJh7WqU/I5pcAL+GSttDk1ZazxhHex53Hl3e1NDLGN1AqqLsYYrYULbObuvb1scx
rr+U4KJ2jyLlkORj2LayWrhBXGtS4ddErDnS1QwP8YdK1L2dLVWeZ1rPw84XZhJN
oMqCjQG+ArzIemKRuGTdkpJqlJOayYuToHmddoCnFd5+jI2F0HzYntyGlhAzqWmn
dOLnueV2e1grui8h4bUm1ez2DYNGjm+aDY/Qx6sxuLm3VE2fKeXzdtt4iSa/Io4T
I30AV4YlfDb4hoDBURTM8h5ihQTb3Vc5kWsZRXQKtiKAY5KbSx163aPakREh2GnB
lzQy6ErKO4ll3d2sV8T13NS1uCNni6gZS1V63M7hBdYYtVHwB32MfLN2sOTZn+TC
YhdYHmyOyr5f6jkOfv8eqk/lfNei2EFdZTyGsUEYC0jFA+37hB1FT6B8dZc3I5Ey
OXOh/W/QNbmq54kEP7JvPfBWrZi+U1Xd7DOSMwdY4BGJkYZlGpkve8Ailfrx5q9Y
HTAz8MFhot/7ak7+THf+VOyDDAcsdHLaknGOdqW3Pk8Ol1aq3fd9WlfvcwdXzimN
Py7UvNZvmsanhW46Bry1gnLr4UuM7NVsqkNSrSOIR2stkFa7hPelPB7piWxS0FGd
wdJnoPrAmIeaxdzpl/r7beQZC0kTC1WJvuBDXq03LLfnEKL8dqGRv6azDjPGNZCE
58cxd/263x0qfct+5unSfa/WZTQt+QYnm1Ys5hk2byzlQz1aih9nbcGnj8CZlYk6
0KSUD2pnR8RTUQ3Zryu2gXPtuwGsLVHfK5aq1CZxIGyQGY3ZRD7p4ZMN5Z7gBKV/
73KZzZz6klh/LAUgYBEy8QKr949FOEKReMUN4o60R6NOEtUQPcqGjvUK1Iy4sLEV
I2KaPRHG2OEZzuYt78vckADF3grZM3QliVDoRcvTHb6FrK5yRxLUfFNZpZ6RGXN5
3SQOSiVeyRWWNd59bCvmv6WNMafC9MIDFRSoou9XD2w7ETmhLl5PqmccITfIxn0m
RoGQfGfPvdxL9fScoc3FQVFSEeMoSzY9/WYhoRG+KCOE5IpMHg/kzngvO+wghelg
bm/ms6bcLvQr6fCWgO1oW4cn5ht4WIz5ahV5T3KVulsofQoC0G99WvonxIT+wwdz
5E39ekIcDSxQG8wZfmJIxPBIwJq9j3R5SFRYXzYyZ80JnFRvwNUijx9JAkxCdskY
s6AuK/H4zXeTLyciO55ODHS66FN0CAx4RpYMRvKk2pWI9L/Fgfmo6yFRPpOCs8Mg
IEI+ybKHiGrRmgt0l30OG/xEVODCufM5mNrmlcI39LNouVGqLDy9eLC6tD5vMWCH
8YnrsOLYcg2xnRBvnApHw801EMY3N3iuBqPVH4o0v/WdNJFaqMdjwVxsty8ceY4x
xO3DWFlHzVCwDdO0i1e8Ri4rDM+scrqdo3aUj5l6fvqeE5YL0e2HIqWvvTLLe/sH
VkE7zrWvtj07MVTXcRQvH2+FwStyHKMmXbtkJXfz3Fxdv4yJ9NjCwSj+SZ7q++pT
oYEpAkuY5w+CiKuiuDeMYAV95Bw5rBtTqeZSSZGPCkdxbxDKF/jhOjyhrB867jiN
9tS/J1YiknPHUPZQoTqvu1k3d7SadCNVhKL/x9lTJWvFA28QbUe70hMtvtZbJ3PR
iUMJWSrgi8ZfxadzagvS0nJP53hdIcOUj22IXX7IVCxAaUaCw6JZ1VYC3oU0wcvs

//pragma protect end_data_block
//pragma protect digest_block
zXfc8cEatlazmwpmzWmr/tv0zhI=
//pragma protect end_digest_block
//pragma protect end_protected

endmodule

