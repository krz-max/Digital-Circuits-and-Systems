//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
p85H7kGz2GZ8ZoMixK3oEEbnS9MbbDAIjQa+Hn5liVhIBbljmT8hfe0DwkcaBv0g
2cZoRIeEVk/MwQMju33WePV+zPt+oPDDJVHRbLETSRjQyk690yPjDe+pFmnc7jDT
c8EfZ/4geOTm2VAXa6NbhcnKi0fogoxTtYqQ6RNtkCoFHZHG/zqkzw==
//pragma protect end_key_block
//pragma protect digest_block
rXeQqolTy9seuUTUWDGq7zF04mc=
//pragma protect end_digest_block
//pragma protect data_block
QZx6bR8xEN/M7ZiNcJSKOOUXWwAmbYZ9/28Zx0t3luRmmtByfM9bJ3WYv5xZ7r3V
Sv8sy5u2/JqXmiWanaz6FXEPPQT3EOZyQCcQfGUbHatZhB/yEO0yyK3nwwihhatd
s0cDNirb3Av6Vc9+XQ/hG8YQltDfLcfKdq30dctSv3zn4bgCnw50to02ZUg3hwJO
8QAOMWRhUObGwASueANk/VTboSj0pal3g2K8e32wsxNW3q/nM5LwRxTBBp5/Konz
3YeH7qDR8lK82f0wk5huCNGTgMz/xLnDgwuf9n1NUbs4SgM+2WOqPA+ijh54Ytqu
wTEViyeIOgC0BFid8DkRd4DTgYNH2LvMJRfSEuGq14i5CZwwuemn7k17AiUpt1cj
AovaRoSxuFz97W8kRwf+7WidBobzANwpCrD7pA6Cr3vWN4QPY8RxGbkqBrEyJmOH
Nt2JG1AqKKz4I2rjb7E449LyZXoKF1epO9M5BjpxX4NhChRSE5senVpET8CcnAwj
2Wxr4bruQE0hourhQjW33AsUvN0u/aOhnmFMTb0hcGwpgZMpbPceEdNVLe75vpjy
jA+KXcII6La90o1EXhJ2tmlF+r6ZGR05IFaWvAikCfVPX+GxDb83u8I8doEzlFfi
hhV+iBawPrzlZpYt2UkZVSRdJKT8278aKw9OOnfzHFz6Yvjwh1eZ8wvIiDayxNnU
wW1Pm0BE7l3Fj454lAjWsaYINkByt3gcoBOKjhSxKvYWEzsia4or0iLscWC4749Q
hsjVS2hoAow+TvQKrLEqYZe/Puo31hA7t9G/AA8Lsw20FMLTyEbxO9z42hSQzAE1
1cyyzzzk6Za9uxO4vNssrBaAKKuKeBf3aVpwf1JZm8gkWZbtccFhtfRHHAy+8ZXN
WKr6ZKF6IsAiPGyjf4n2vTaR7g0DnKL0wtkpH+4quXs7F+oIiNm75CxI1dbVofoL
sS2PFR5V0M9itgf3J1ydYd7foX829yjwMc3snfBENXcbegFDPIuXEGRBkp0TJxOK
NpIQe2irwj37xs1IiG1JWHSiVbcN/St3RZ3BQdYB8HD862YI54P6pqsHvn0xFt+Y
TicnVhAwxuzPKb7ZJ7Fn5jYQcUKXXqGao/kMSIKBRq8aovryykJqe7zOW7rACERQ
f3VWXmb0ZgI6QMdO7p/IakVDASdkI0ImrjX+JhblOrTPNKdzEbAdUfjDkL06e9Hy
I/XzWw+cx5+3cQxW5JhYAn0k9g8Otvj+2rXEiXwfi9j91PAv8Urh9z4gxFZ5QR25
oX8Bk8wcrP/WjaZjYrR1rvpziQHy7gKk+m3dqsOF5ok/prNLLOSZX9a0FzS2MDMW
loAemItDGGI5MDwVDUEnD1nDXcciE5sgm1BqPxPzj0Y+X2PHHOgTjhy+2rmgX5jm
lfFBfcn1hwBhYmptUyiANSGpogfqYE2fR+81xSvNwOu2DDOieV4Ro79PTjO3/kGx
GT7xs9i0FUuAjpFACRwBfbK6+iOhlD/n062yP46uTCkeR4+DOL9eOKCdO8nc+AZG
WBDMZfJ55Q5IAxKcVTRPFrl6gOclIafTa09Yqhq7SD24vq90PoHOJB/TbauT+AHl
1rld1Ife87aBgD65cVWD+yp7oITe6yXPL1UUaYa6/7wKuHrglBeZz65cWtE2BzP1
yeoEimaVKaYZxSfprzqxTZ/BQhQ43f1eObR+GqpTKln146jBRh/QdvEX0HQOT4my
PzbCxOyrSrmOuoqeGixiF0fXO7+xEZAxeu0t7LBAQf6TPDBpcuFP/AfhaQNzUQ19
xog3yB8hxAz+C9wqDhIeKCAFIsYvqA1blbERN6bNvx2tO9RV+O6R4o9X7sP3QDtU
TnAh0qVEdXC1VUIqCedvREoL83paj10d4ENC5GECaFWdqNEbStt5BUvhPs0VlQFd
hdCRu5eZutHbsxJa/gs9ts2hem7sell8GKpMC5OC8b8G8opCHhHUpF8AbKIWvR7s
EPeASutE/rUISBZck2gJ7YXQ8dfXbKGBKG3AUdyyBecSgipseP/WuwlcjkZRivly
maD0t5rSsKJ50EFvrWLMLNL62lDnLmykDylOkSRMpl5ibCKG5JWL5z5JOSL0DMyS
WR/CTO0mN3Tv/ni+7Hj5VWgG7WSeic0bYS2aU4x9YzeH9v/1XxYgZy3WlbY2P0s+
tVAIAO+pm3UgeVmFYVrbMcF16knBoQkXioy/1e83UQIrt7b5KhT2M4gOMaa7tLHz
NYonI/mwUt8qP9eJxQgAJKgrfuZ8pDbqBa7Yp4sxf1t+BZY5igOBYy9s5EI7Q/VV
O6DI92JBqVkhN89Ap4QaPM1QtvnRJr3QHDMm9wBECERAIn7HIrAjOqrVd8nvgSk9
VWMS+kTT5gQKAoZGN+XZ6jDTwWkX6+nQQ7FmmjexoAlZGYHEtISS2/yMFnfINBqO
dcG5GwQZ6c920o7YJ0Q1ASqcddBVvfSdQ/uoCr26mCnOmzQd6Nrd7A4rNuWYxC0Z
HOU/rmTUeKiYbBi+hIVZ05bzxP7b55XsqdqWiBQpOmuU76X+iIg6nOuWkWTfcgKv
JY0y9ikC4xA0VAg4aXDuWEtW5DyYgfyTk8hnDguQlj9kg+6pfJZTgDAwjA6q8aYQ
aDTQOug+y+oMIO0C/KS+p8P+r5ifgDmfnd4WsVxWypzWDg+5Wg5+Ft7qi4TaPzVv
naBrFEScC2U3OSOm2abBmj1fvDkKY5R9+UD0xn+fGzzfI1KKbYu2XATT4VF+Qke2
RSIyypsS+KGa1dW7c8jSWF5fCnIUW4QEOCRyHE8TkzxmZnE9diXdQ39cwK0qGdNp
vmo4SOu8i+ttOQe13iVHuaxIjFBdDuCAESdr749T7G78noHZ5QeqET1VQ83ASd/2
SMuyfp86H8iwndw4dF2nJrPzBnNkcN5F7ayCe4nkLlyQJS7O+Y07pVX8rWoipzlw
ckO2BNwfdYxwkeAxHTbIxk5dzOWhOkAGhG5H8xupIw6OMbyPEeoKMWSB9DAaBna/
Dzm14kJLfg3uQidT4K5sxzXr7+QBiHZQ3VI2dqpK+eium8Nti3m6VlKbFvkRYIo5
ts/0qgv/JFPAC2RE98Yd9huQRuYUVB1wy2pH/9GOGgaUbJAYAOkxMyr8wTzanrGM
RMyfdYIznLBIVQwAMXYFk0IoC38H2VlDyrYOfd0//nbLM04oCTiH/qnFWLHKPYQi
dJZ5x/SIq3HRcz8FCMkehKsuuPDs0V0w/MQ7wRA3tuWquhFIQpRkB3TRwp4bA4Bh
B62vI5DaoTQJTv5892I18Hon3TvIhwrOEf9LY/+3zPiwFFfIhyeYygVLmJLSgdHF
xnWIg+3J7hKYnArJDotHi2/OXEUpgrJMJNX6f6s4px5mTPlqZuk13K9jH/5KcvnC
wFVCXB67k2GkVCRPmXuBUTisIoHqqElpk2OS7ND+GzInEs/lrecVSEBKSaEgOJKt
RtplA8VG8WIfClj3LoiAeZqDquLhDfnmIIDhW/FYGQeOgXbRpkB93IKjMOaWRyUf
wzbNZPguUqWPrU5itTvWV4+xwIZxje+B5VFZo8PhOZSu9Op3o30zKWpm8bIqSP0N
ikaeTrdH1fF2EfsJG1ztlUWnSNSFUN+7llMM+yUWKStGqHRgJ9CdY9e1sNMe5+9T
3UIs8TJuehx+jbpEPeOQ923rU0mO+4SqDM5R+Anja3fbWjDaVjC+U99xMFEGkYZ0
wGLac6l1B6wXjMp9NiP+gTuWjEdcsEOHLNgH5fNPOIg2A8i4STv3lrrUALSbAMx2
/pnvk2CnK36pG4FFWar/jbrJXRqV99SGI01WI6OVcAX+YSibqiPaXNUC9CF5KFvo
HsYnvzBpfSzZKNT0ZwBRQBXONjJYrjyudtQYNacOyb/Iq4pB09prUuLcyBrczCQ9
i2aGUTtSNKfanfLOjUl/kHzSzPTds/IHX+USUjsNAP35iiD8L37u/wNSY3lH+X3V
Jl5JZ4cxF9UPIzkklpKWGKQY5MLJ3Ar0UwawfKD1XPxLQLz90EgCYnNK2oLCrk34
dBe8lGgf+VzepZK0R/3LdVUshzIPuqGAvVsH/LS4UIRnlNjA8Tr4OyGYaM3gxV7w
vnzax/zOyHuqGxKfKcRo0fvC8R0TBuI22PrhQZbamfrDWwpRD7Jq1Pit2FNz8Qsg
JaKtYqZkptuTW3ES0A52Ksl9sxy9gfMG39skmzKVhmoV6DMwP91oYbe8pzMPT6Uo
nOXs5urv7Gn3D7+U45zs0rl4VuXokpmhHIjHCTYKTSbmkdYd+zT/CBFSKsHJG9SQ
xgx0MfaEVPmr2llau6EqJmU0MeK4YCGs92bCrgqi+KGeSCXhPDuFO5thJ4/Mzf5p
WCpk1pv5qrJ8ai/+RrfBGozDZPhRy/wUyl8fBXqIJYezVj7ENYaBBLJ8wUdjzzuU
aSig4Pw7Hcq2a/ZAVry4tkvJ/b/Kn5R0rRfYujXLKz8RgAgWU6u1kuV9F3U2RqU4
PDvQ+hULqlhB+OCks+JqxuROn/aeQlrTk6XQNKlz8q7KQ/DIruwCTTNta/SJHuvs
MCw0fQzMZSa+VRb+dsRrbclnZUm3WX6/iM202qSr0ZNdJlET7meSxc3tfIkqMjjx
IOmrC6mr/Z61CeHI50/SMroArMLHOvwv5T5+Aj/BtYHAhb1HakhARDKFd/ZUICqC
l00wUPY5h+3aOdebpUrriMT/NCHk8apSAEBGAYPt1or4VJOqGkjQJbbcQu2+plfc
O5YHA8uDnZiJSfA9qjCPM8qzeYuJrtIY3sdz+Y4QeFT/A+h+EMPZZBEn2+KdSeSm
9d45cyhzpnUnd8awHv3/CxepbELcWVqsyIz1gzfvtx69ciW1RKQa6msKzoT2Bjy7
SREQ+mAtvNRCe/7M833LES6glPPlUlfZkBHmck14XXsd6QwEn8Q2hY6dysPf/LEF
4nQyTrJbkQ9KuYW2Jj1xQvlrFBIkqR99nndxhX+qSDfyv5mf5zXhSVHBPzBpHfQV
rq2Zq8m5LmVfOpu90DHlIzsRfbsMGgZE197RaIFMUKhZIT+jjjKRZgCFQcznfa7q
fhDu1AgpyQV1atFYd/6dS0Yol682hbUGCDuxtQXB6zIbRfjNbaeuqyfX3ZIjAvTa
mE0CWD2EhGW/Lf5EiaqXhhJ2j33AHZkE1o7KgO+4hlispc9KtvzyqAkVXKGe4uVU
FhjRISEGgDvj1zBtp+P1bFtaANE53IihNuuFgT3GU2z2yBsXh6qggkoJMsoIPHOR
j7LK1klybGZZUCjwWMk8NPbWY6pt5EogA1XiMKepXNI8Uw1fhrHcqneo2PpE31nh
DJC8aFauFz42StiCaAWQZENgjFGR0Mc4MQuIFGAtatQvXg4LLResDznZwkL03NPm
fIeccy/g5ATcYUWwHpjLinnhKVUqjdbemHrCdfMfzNdVDiK7RavpmEh5stQbMx+x
OqPh0t1V9IBXg0NFLttp9gOB+mHRWFnebZ9CaI7MigjO0AKpczHSJT36kXInFr9J
AD9Q7yQ9Y+kTYfIv7n7/8ptMBFjAaEsrSgUkdn3qIqWEnkaK7k5VkzE4IEgnNhCZ
4aUvjTnKth9BuPjoGB/7wn6krFqw2Jie3jn/QGqrqT+sLv+7zyhwLVACGrdXA7ep
g3FTxUdeyPMEvAR17sHMsFIdaNrEVy+vPo/LI7NMXAAsIvnEYl/qrPzLVkiLg5RS
BZCecM3nhiXvXr0tip+J7Knb4L1bHvMzmQjRhaQXIYmDhR/iX1ruHZWL0YkRYQTj
mDUz06xplr/TQ20G0l2HEYyDCwaj2AIk/KuHsJW1GZvXr67uFrHAnJq1pa3SI2Uu
iATxt8ZPnlTChlzxY8IsWVhyDzGQopCBRI3x29Skjc5WSWLnBEgdTW4/jRUNOaMn
f+C5ZJYiQln7jQVqaHkm/B0LK3wDKSlkXcurQUxYavfg1IJu3igXk//d80qYXQ7N
y6xvgk9KbGeOZFMGIrWG4YViZTnyW2Co3cXEIfhbawR9YU8eSJ/MqYcjakybuxzL
O/nDqDtWn/nl1AID0+IIQ1k9okjnJQbURz1EWb//3JIAfwmqzowxGH/46DB5StFY
imHWocJXF8rN3EZ5jdwjqA6taluTXhWQLCLhUgrAkuMUYKLuRlIhHxV7cWgUbbRr
eUjppwj3C+gHqG4Se1rNcSl+AyDOI/DBMmHwgVieYbC3hzhl1PjVOGDOEw3H6nj/
lyMeP1Uc/hhD7yRZgjzNTNZMXVA8fNYXspIyLKjuuPFD/bskU8fesCqiraPCUO2a
uIYJvwxXcbP/W4KQ9q6ayr/MeR/+LNf6MDGJ/Z0/sK+VZIiL87BlhGJ9AhEyPzJt
SY4Q3XeWlDtXhRck6Eds1e/HvuWU20LTk8tdUwvUhjEzBtVtr2ICbR4EYM+BzUxE
cgh7Astw02fGAO/z7YjD9Ogvsnf6bgrh5Eytr0p6Aid5AQ0bmUbrYDFJP8fFGjoG
gmzyN2LWETQ7tJIkVqVziNb8HdAdW38mBfvnt2oyhThca/7DcGrF7D/HXQn7VZiH
nStJBLFJgqssYX0Xhq8Ofn7tFgrxW42R8FpHrlEYs7OIiqhT0CPd0OX3KFStdnPC
FE0OzRgAHDQThaMvzJ+cMv6UNqUXn3ZSo1T0Yk3FFVzkNrwhCpHjx4JqAW6Q48QU
egOmRcl+GYli5AvCJV55u90urVcATehyeTFQ0sgX4ds1apmEHMG4BfHSFuoUfxmq
5GGjbO5vHB+HMBA+zYlDKBTFxF1Xgr/SRwiqWnSe4aBWgDgAvrOH/lAnu55y6Qg8
HSeqk0qrymH5+2HG18+mEHJaWfU9WO4+VLOSHMKMfs6KDsdOjJwclOZQ7hoXCrL2
xgg4BvRp222fp8ffQW/p9MLkVtXq2yixvJf/Ly1bbqOJhbM5bID6QvBIZDG9jrkw
esGQdAZXZLFkAzVQm5E0KcTuOCgzllXBLPcIhwKt+HyqAFLK8omx7Qph6dB2xipo
Vm/bnR6ywbAzCsAOpfjuv1OOphAs7+P575ehTbyOwXkfoJPHQZMDi4YISBpa/6sl
PdNIF0ciyURKYvLCgcD0in2Pxx4DdL+ghWgptynhO8V++c/Sq9R3O3OqtiiV4zti
lMTvVd51NWvjrF3vITd713PXn6ChYuEvrrawE4s4VwfVzmZh7kPkFQ+vrwwtEIZc
KmvkbZS/lKJAz6vubfRyo1JW6716Xi/IfoGTtDUereD4BdKic38gTLvcuxSHFl/a
rxCyYz4WIJN+WQVl2Ke9XT5Qf/sxpLIzZJENYUQGPhuFVd9RFuOJB5UH0EE2ZQ49
1/8YwynY9VKalTrBIcCtUyhn2rh1bus0vWgT8mxkTlE=
//pragma protect end_data_block
//pragma protect digest_block
pTJBYF5cXSAYOM5KoLGWMB2pRZE=
//pragma protect end_digest_block
//pragma protect end_protected
