//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
SaCaTWQEl01Wq1fXmhL0ALOOTGnwc20xdfi3PvsNuWKkmeOZpGFDpVhfHu/VwU7R
E3axCAZHPihKpHIZKxCVlNHjk0k4wlY8m76aQgNaihlxwQMR+lygDYe9zhocaEl2
i1ZszgFGWiqk/bYYuIr3WzdN7f+o2kT2WXCIxCrQyOpap27S9onbXw==
//pragma protect end_key_block
//pragma protect digest_block
foK++m+2+qWzraGLMs5QIXHzVaU=
//pragma protect end_digest_block
//pragma protect data_block
s9+67/D16GnATH5F2Lu0BLkPn/7DoM+ESaDU3J9Y1EoLj1IEMMQm1N8hirRPwOsD
7zudviSKfl6RwNXGn+9KNNNqwCJfponWDjIRbuA0Q5GD5UPK9EdXG28zzYNXqwDv
lrwxWzpKh4s2W5ZMvEHxW4bs5nqgy6eeDjI/XUeu1+AbCMb9gDXhTOfmsvFV4tpp
6IQv0473JrJyn2k3kZpx8iRN5+g1hWL4DOQp/L++nccyY83S2xCVlKUWlDiPrZl+
/dzpGam3EIa9YgZ59dmu0DVcKGKOCwRMWE4rpNf7Emsg/hnyD+wfcQmgPmA/XX3w
vka5miGMo53IO7KFImmxMqoSScrqEWZPZwzbKO80q4U4YHY96uM2pDGo94OJcUah
1q92sEJbWRz+ycEMGB6o0U8gQRoEEMH33T+xVG31TfrskRFXibizV1QHimf3WqvG
P+TFXIdYbYq/qiqjKDirqvUMqiEOoV6l/R7XDS86DP5GIbgiESlwKH8YXd+x8LW7
uSzOTBHkAYvp36qCDRnomC57MudzbIPHXWyqce9x9jbpEi1V4nrjLeo92rVnflDy
QN7Ad4oaerScFdv1ahatoGumz9jqjncML5TdSYjeAXaUw4eurpuj7QX5/0Z1iLiC
jPIJOGjBxGD8uUiZ2WfeXFgdPi/kPpN8ONXbf6nyBDJLwWnNeZjm0HOuUP+ZTLqX
cAAHLcuXrxwLGYjRF4dg8NJLXoNkCsjwTfqY1rBRo2xaLelEiLWCvTmIvrrQjsAM
SfnBhziHwDZhcz2GvgqPpfKlinp5d8EU1B3L7kvoYbbqINeMCK7Zlyyo8i/x19SO
eJCvU4yhdRHG0dLS2kA3kh+6TV/bRHV1iLysnin1Bcop+Pwbn8X2xLMxWPedLYr5
DPzGq/s0QLGmdTFb0rOcQ75NndBLfFnIr+SPVPUTMljsYouJb9tlY8XJfXdVYjr+
iK2uvY1rzu1MvaX8OwwGU7j2mIcsZI18xndGE6utYlosL6axfKrQ+BQGBSb1GHHJ
suJM399exg4rzXCr8d/1FCTTc7//n/05BjRjBYvf2YRHUpnMhZ6hJLxm5LMqXSyY
ATcY8GDZSV2ioUu20WDQop8YVP4W1wkOoyU2IXr/Bdfyr8Us5AlVizppuJ53aATX
8cpGizvlzMiwxtCmMHKmz+RjClY9uS4AyuX6Hew7njneizeLrWk1hgh9ATwnVrEy
4yzDvEu3XQJT6t6uF3JTXmAfuLRt60+i6GCQfd/fjeEm6JMc3SXIIM+DONxv9t/E
ySlfGyB+bLZsAYMXoRBujCySgMVNtoWHoIW03TnrZfLPjX5nN2ubKGJiYUiemYD2
u1ZmWoaStLtzvBvNvOk/WAEJu/074V7S/lsxBpFgeKV+z+V6CnQ+E56t/IEv2PBM
BpB+/d5w6MjlOPaA5QGA8fAlOxBewGKuS+shgp79y6cg1OFbYbwNGwPHdg1/X7q1
2/1yOyZMAZX5KU3EIgXPMNky4TlO6lzAPtpBRpiLPPQq10QdibA6qudawLT0kLq9
7zo7E8RFSMthydLROVcyuIihg6JLJ0LAwZQ074/Y/RY5NJoaBbqvtrUuzPby44hz
UGi6JFIGC7VKxbwrDnyXKg+5Fi78TvBsKcBiXvevYIU/nwdssmNHAsDsoKL70I2z
IldUd57QKFmmLY7Bpl5iWub3gIeMDpD4C74x4yHsIvhFTmzQPB7G59rk8v/PKBX3
S3gXf1DXH4VCGMdMH9A+9knVtN7YjiPpFt6pwBoTRdC5TSOgFWXqSxuV7N3leEzH
3R5HkCbP4s22g1KajHUAucPnsV1OtHANuDi7H3XHnw1ld9Ujm6KhyqY9iAJ7dJNF
lU9gugjG5aSPZpOn/wvQPbSn9Hxya4iGYLYAwdWYu7e8YVwLTK4Ni4T6TiKfPPsx
LY1UXDQzZiUpJ6uOVHS5TaHzmvwhlMr0OYJA93KdHxL0IMY6IgNJHNXcaYjD5Pw1
z3btogH4HA7MhG1mlJhyF1848acU5+bP+9WOEs5JQFG/7JOizxH/BZRi5jTJ6yJy
8Ij6T8ETfYDvkxz8loKj19KjqT5azf2aiI1N1ytDWcMUbEOskZFZ3vTrSWjOVLAp
0ouICrXNfnjf83P2tyWNlcNDOO45c/s6QcfVARrrYkSeb6AkBWiPFPlrBFg9Pxpv
Ej4uQcikzzSGf3sA0+mgSgDd3AOHDl5P7qFMzDBT4ujHzwzFCv2ouOVrV3nktrSS
D0fIu1pN6PJ9PRHEB455HM4UO4kwLsaZyzE1eRGkJIZFOgDOPlrspxq3Z4rdMEXr
BV3JAIbtfgm4ja5sFf81UATzioj/TS7SPX/hFBbIKYzpf+3sD+gBbvi7BmNUDDL9
T4VUj0aYYyAyVjR9/w0kw6cgrsmzqfuE0Uy8YZq3yk5hGNsDp6r9TbRTHXroCEeF
XLf5E4kZj+2D07N3FfR2Gk5HJqsvVtZ3AjkkPAO2oY65PS9gbc1BMtCc1qrN3oAE
b3y3kUAN7YrwShB3ZpCTV2Fct0Fu5fILB8XlCTHsvIFxQCoF3GBLzVb5nxxsJijz
Rg5P0lY9h/o0DhZBE9W4JO/o9fi1ixOGS9n5ZRjP3WGSvAIc8EvczMCuIfmchFRr
825vz9c6Um5H7IQvNRajMAd3X/quF50xVVBXk1NzpMn3+i8V02xrsRyPyXEwEVXK
6RxPGdcGB/CyrfuYP/4VQ5IITKYDhh6Jj5HKrtRBy8YFDSYuB8OEu50ns1GoYsWW
EOLl4PdRervNLEzLVAerJD55OnsokEemr2NEEouBpHP8z9ngM3QFVa1wyFthtsyD
BJT06WOhZJrEtLD66bzBT1FHODt1pemjGO8TEx2OzxmFAEAGyC08386EcVy3MYEu
Hdewau+TJBtcgSws/rnyzgZEFeg6C82heqP/z/3dbsOsRGB6sL8hvVPaHjuqUSrL
n5q7zQ3LOfG/opSamPrGnmJ+M4cogzzg+Q7Q9ZxhOg5C5zfS3lEmqNnN/uIWZ5eG
cpKUX5QfABf/IkobVgXVgflNj/0VKykhc3jEA6YNjK9pRtCMbNNf/kyC01J0AUZP
uKBKrayjnXwu7lJDp5q/oC8HD4rqv7Ab3vkjTriNYFyKdzq1GS3DldJ35dBFd2MW
Hmio1wKmkW1i/9QKfd3UQM+nSlm8LtNPJsfqMu7ncPlb6uZLE5zPqbb3Uy0J5TbK
Ohr8heFdpJBkaishg2zpopZbaRsidz745kI4vznHCCz3+e2cC3ovsqYim/q4u/9L
seW0J/mJkOPREOjHw4L45EFd8nGzVvgiNbTi6FMIBbxIU0vJ5kul31chFMAdX84/
z+qNMBeHdaVza3JJyx2hFzXGIAKxdbrDqOJ2OQRkPnwunV1I4zSzdw5DPewhMYwV
b7q5EncxlUvx9TJLT9k7PAXopFL7umf8e1TAzJz3Hzy72gyZgWGtFJR5GXPnr5cF
JKikhPVcyCJ/t+bzyxnpot4Od5EW/38qUfxo/Vg2vOKnQgYrx0NUSQxLj2u7h3s9
ywXr7qZWEFgTRi3YBPrP7bIXFZib3kfxAhW+I/9/00usLq2FUaEhsZYs+9mUA/ue
mb6jnyIPKM5qAnbSbM7yOcRjBTWJg6vtrIWrozJDqoSr/nGZhPe95lHGCocjxt0R
H2wcasTtCUcbnY6DyUs7QGw8nHr+vpSQimAJ5UWBEkFdzj6GEmmTKS0IGzlRijS/
UP3g6cvIIf/DSm0PMYecidEGtSX7T4DQ2ph+wCSY3EGVc81vfKRpGbqmG9UurILB
mRB9uFROyEhkrsUDFMTf52zpzsiAHkd57DPry1hT3eJ6eHBu6P+zQIHc7UR6Q4qF
rHyu1WclQcsPbGdy8YghPwJ5LqQaRyX0GimKW9nSuKfc49nXzBv077g1QrZrgk+c
o71B38jmgE0/mjfE8NABqbFiY+LOfOlt6iPDi/aoryRN38MftII+AfGVpdATpRjY
lQfsAtgv6dN37UoyXhYP0VaY2a6bgbq0ZEJH9QJ20enifVsWK9PirZ9AxqBnbJb7
aVjU+fx+CSf3XhrMX5J5Zb6gV4ZisUvbTz4UZLkvX+uj4xQcKOSfqJ0ftQHmPn6/
WnjUFTvcIhCwuMPYHvcOvw4nHEe6+5XDE8LveAeHP9XuYvmukdjC0jMMSKr42Mo3
E2r0ZKJAWxuw3/ssMjhufxj5j3PcDUtm5YNqJKqKi/OBhnKUkipCCpFR2ncTGK6t
EwHvQtzdoBrHCugVcK82yOsqyVZfzsRiUuS8fFtZjxv9FITYFRfJ3rWQeDGAiSYJ
tcCjxU6L3/rFlWR+CtFs+CFM0FXPOnBolIyoLTw/n3wDuTfHG8Kg0+9mnsyiius2
Jsed7mt7xSBcs+Yt7AcaK6W4q8WxHdVOJjCy05Y8841bRrDP1xiesATriv2XQxKL
K67BjZgCzRaHOYqd0x68sg4Kd0y4luaSjz5ukqTKU0KOaYxWdsphqWL18qbQxHKV
x+RZlbsSEwgFL50KQpkQN3CACljK587I20UYmA51kZLtVJa4o51Rc1mo0ssH1dSz
T6rsoHXEE9j2ztwsdwEn5GquKsjXK0CfFlfn5XpQ+g6bpjEDd9gTfqZRuXorF1G7
nadhG49ChoYVUPKVXOVnmKtiIQUfJCaMvU1auiw/CO+fxXTxZFedCM3RpXTnXlP4
bwwLiBFNwNwIJifS5MTi5hbWDav8ew09l84rvWm/D6m+TLxIMiRr/BEABWEn6MCz
TV38gQ6zD6cPNyt480cuRxoyBcY/LClOjoOpdHg75lP44uojXaNweLHpgJX99vxc
qgyZDFGvfdXdzWh6E9QxIujC9zChhASSYe9HcyWCymyb9j4D48qVWw9ttNvb8rMY
ZDTTpfLxPOMWRVk9TcOTN6HXrXVJdUE+wOsqZTmlE1AdyajAmtH6lIVqueoIG2lv
ALmE9i9yRD8vcrBSUumxDMUWOXmqZ1fO1iNPgmXFMuZYAnAhMuSN/HxI4cthPLnh
Kx37nf3mJnSGhLtO98nqwr9LtTUJpE2mDvD7ibeXunTqBzLtygE0PzWOmTVpyGN4
ke0gU4wh66mj6wxNAD9CxLo6kz6jy0f8l7uPAobHnsxSWx0xh9l6uwEfXvGdk57z
icA+7UQvGpKbUEW3sdzRiBGxwUxAen6+uagqI7wElSQZIV8JAdF8BhOKWAfDb3Zp
8SZX03AwpNVq19Mozp/Q+eUJ1BCEaRs1Z2ukHrJr27KxFBNLNNYTu6+uACKmD1Cl
vJFtE4P5R1ZKaCEyz//+aqv6fcsWTjyN9Px6E6KN8l7P3KnA7bf4Rpadtnpnv/4y
p/fSbGojMJBAe0WhQoLJA5GZbXfldDGobFMxEDd40f9bQKmBTWVsaMmhBAgNBQYF
0mwi0YBA3LjX+PZYFDkGd8dPoNIY8NNQKmLVpybgoFlBi17RbVqxxmI4yVQ43ngn
sIT9DT44/3cVDQaNi7VTXKjvyb6rql2u+JU58O/snTZTp1u5RktSbDdxZ2o/zsYr
tcACnevb87hEuUsshW/WTeo2tEyNRG1P8uibXuR7MuYcPtCs9xePY3BVNWtEXqNg
hGKPh48ckj1H5Nn6aHRtz02kLUCWybMEXDxFPNeA7Baa+JJGhvSYW5RzMxxOWZVo
rtljWPTEFAvvd7ciRqGyGJL2vqfsE+jCgNMrhbUOhUWzfoob2vzs4B7RPCdtRw+A
J/9eNo8aoHOCRKlOJgcm8dTqzay0yEB2X3JQdJ8f5EWYk8qkMHt+TZxrGHYY8quN
f/TotPMQmsTeUs127C42z09Rbd/HZFq9vzvPoLO3zR1EG2dZb7WW6nrshsIaETA0
Y/eFOaBjr82VBU4e3ndCbFtai1EVVavyncjCWXSHjpMvnvbN33KuXW6RDhlVBtHS
LB1uJEv7DMYQe++xHbgCZWOqsXfzRkc9XgoBb2UP374ESsUod5c8pHOYr9LdV+RR
4FEPQnJxMeBdqjW0S0yH9YjQQb9A8SMcW+yubsa6pPOXUqCxHddPLBaT3gfcxiek
KoEnUr47+8tsFa6q1cBXaos59j2Wo2iivEeoqG3gDvA2d6RarfTSAjb1+dmLfUYi
KaRPzmFzVqjbblwKIpQaVDqTq/YMLJIX/h31AlsbZF9/grAmzooSGSbxJqqjbSP0
/X8LnPZ4GzDokerr2LVd8LWoCBMwFbEI1exqi2VFda7ALCHXTgaoev/ZD/3wzk6T
zNg616xj6A7WqVTXBU61ZwCM+Tks41LFPtvwLp6JDzT1kw21Gs8xkfJrIIniQVYa
TzHvo+ObFi+nhjDwRIQTKHchByVsmu7pm9fRu3iXI43kW9Q8pHG/FqSjC/24j0gW
ucts2yjHIVSHrPIFn5xw9WRCJF468nbQtZQf1VrRDRErlEahy/UPtVGTKXMkUJln
0i8iD7Leied9ohK4En+nw6hQSF95qtU62rR00c+d/U1YKAZYBVD/yJFRR8sv2KDv
XeewN7hnFVfYOWkmLqUoksDQyqx9grLOmwpAJdYlbEFxsoLUbnOI1Hvq9mW4MR41
lIrH5LNsl3KMGTJPhDF03m+K55T68N/CSU50IWO5Swqj8ESjmShUxVuU0klgtIla
H1g0BMyPLz6Oe/wZ3cs6TMB/ulPjPbytkWiqnTkOZtdbfUKnrm9/Xdf/cv24wxqH
8sz0XFZvDJTRbZQahKCz9nSoi4R1PGZ2xvovnlQt5VXlRcQIZFvBzxWKQgSrjh0s
zirEPGKIcZQrMvaN0zxBcX7YWP3NyVCMqKd2W3VitlpyhjzzIlf8RVyt+RIFcqW0
zdy+J1miDY9rJHAD16buk6YRfmGizws/FUMpmQdZHfeg/Db7qB3jb0vhr4ySSxFB
rcHLBAjgY8zOPCYfHWYZFjqKvyDoHXV5HSLwKFqGjKpPztjqYYeFCf409KQkjiQQ
Z2VOljOB2UscUEazWS3HCeee1fi0GUS8AYbvubJcEg4uRN08eOB449r56TwL7lfy
joM/NCc57NYR3aWsQQQe8mT8CeJyFqL5idvDWqjIwclA9vokTiyKI+K0QgJLnxa6
fh6N7tNr9nz/3uCyQWvvUYkf+gb8GouNpZE1JmzBCYUZPz00By4yOYowtvmimlVr
NuCSUYpKcjTQuxcZNNJIgwqB9Zw7OCx98+8wi2Pkh4+/pjYA7EA62Gr+gOXv7uB7
DDh3u0LhMSMuG4lJyHRz/iNRLYPo7p0dkX6cm0fOBKzAHU63oBsCW5FU9UXxoDNA
PDw8Bz2D30j2Evkwh8NYYX5RyOmv8ga+XJxbU1yS2hMWaBB/8V3Oad2FsPMZhUj9
jfyR3EB7dLcK42l4iiR4doyOKtNyA8edQ+50WPRUsXT6JSCCCmJW/I0mMOl4oIZO
48MXwmtgczeap9LdT+uPEHCHWncUeBwYAP2dmfdJsbaF6ZjGs9EPtJQujRGhZJjl
nbrIQldhpNBX7Knp1YpLkplPiXB4rOOzQ/N58VJKXBiwMWZ1QIZZACSf8UiQzUTk
Cr/AAXahWrjMdjmt59rfO/w/8oO4z4vD4lnsFJCz0hBG9W9QaE/+lxUWh8DfeZVI
dQjDCaZFMmlgVjQbzCESEOyW4zEh2L9dtx/IkfKrFlGMQnT8Y7amPnzUS4M9ySH9
MBpJFekH/U1lasw7lQh9cYvsX/7Xvde9xz5cVhPXY7aynEmy0jyCngbxGvNBlFh7
RNttieSIwyJeGlX6MRzDdq6wu9Ep9k7ptl8WfZOn7a9LSbLLySRQwtsOuUW2bQqi
2SzkXeTvArjJlzN/CZiV2jCfKpY/Sg7yKUp0g9/vjYpYpmXKjU1V+wd9MWwlANBI
gro8SKwR/UcA+xzy10V+3n+r+jlOav+uR0ZKam5rEYUMhyTT2l9tQqSaGTOI84Gi
Ug0NBK0VSJpS/q73bakQVByBA7H5dAXATXVFXr13hgdZBInXmFD3DYff4STwyJJl
gRykKakWZU1kKRYjmltNuPSnAO0OPuikGp7VEclwHxnlmkRi9XI4lCzyKjqaqqVX
B7fHiOGP7osXQCoCvkpB2DBbyYMJfNQGuMEwO8a2WrgK/0Uy4Owkq5n7fs2IrCGQ
JpABZisH8ovmAx3xMnd3lVvQu+f9k2klDvVLSKTD6/QnsOdo/V+qWew/fUYZPHCR
Sq1Rc1Wjc3IGF2LdsfCQ1etvfi7fDhVlG8Xd/T3QMQkRVlzAn0Y4i4Cji/bZkhRR
sZh0lbh0AdZ8ZXE2VzwICqde4a5RXiZwwmfNpEh0QRm+QeQj0YLEkRUI1E2+lTzr
TdNkZYhQVr0KMSirRnvZ8YqPMZcFYSc3M+AeiFMDwOi9VqQJYRZMUQ6s8ZYVvLBy
9V3Rol2V1OKtFKi74zJAqWMRy44UGOmtYbqzBUEM8Kad03HNigSdTUaEd2IBQHLN
jXOpAA1vgfIjmbMySJ0f2DcN4exARAFq2Yel+AL6dtAZ5xU4tJVT039fM6lKCWG9
3qB7g8vPMJ5qlvSMU8chxmhhZ6aPWIlkcV9hueBGw3QO4Vh5hrnDeA0CWWYCFPcF
KQMPbTuFo8mZp8RlABkPBo4UTlNQwIiCRr8g7SWdymjLrJdvyxjtasNf8NM/jVng
Nv7jBlH4ZIo2F2o/CvTBsL6LS0MLIiRyGodYEXCoN68U6pEgfwp0cki5MPr4uNoY
U2myW8h9HAh/+aY/QIdn/nvgFCKziVYhsas3qGBT+4LALAfahyDtWNtlLCbDh4kk
jbvtzjZPmOIpdnnURYChiHHhXM778aznFCEvnvu6KoVQNLf6AhJ8ZcVLvY5rl1Sm
m9Y0vU3FsCP8tcq1LDf1xsswG0oFVTB6S4EltHpVfvC0yKwFCE7o+ZYPjfpN8u2A
WoNnRkbdhLtGl5HHUd8GQWPM5yf0Mtk/HwTwpESxKiY/1swKiTHoPO3Pct7dRxT/
mEjZeHJ2slIWNSCZnJGZq4s9qx60v+grnU9yzLu7R+8bd7fAk/nsMT0If6HbU0Hc
hSaSUELlQW9pCiiSUv59lRk6qm/7REBecEkVG1zd6oPyCycunUeOHNTtlDKFGQ5a
QZAqJj+GTsAx0U9IUtEzSdVjnZFhl1TDZyMQB8FVJS/S5rOqT5hApsTfc5qDeAJV
MSXjnBzKWskY3Ux/NqjlK7YQGgL5xuYzCbtHS6/ZTWODT4dVPbwxSrOcEn5gGkis
UtiOgZkeTM1You2eDC8EebN2iB2shgo6yHGY2CL/2YM+72avJV2p6hSx+NTKOE4o
R/2yQhZaLYymp2+wctDxZKkjcnkHIWep5VAlnB4oUIb01NMJ1205G+akicNi8v1P
weUDP+KyNlmDZfYQIbh1S839jjs78W7LCE8oqZoEfqdyLLbKike9OgRSBFLJOeYN
SIOaGjGWR+PE/7NGEFCUMvUS1QMt1M0QA0I+dDlUyaWJ+E7IeT96zmz3HbondbYx
g1GyNjWAwJe7D6G1R5KcV+XwbeD0iKYciUXfYXbWm+OxMAnbPwdgylo67B+9m+WJ
mTEXoQvFo+RsL5G0/y7EIdIfCIELlghIAYHq5mcvVyVCd1h3p5lf3liimWiCqKgd
hNS/ey+TlVFVAQiATzzzEw/GNSaTUXiEPg98BLTngv05aG0KCgqFuXRxoGbBGE4D
jIsCmieUFpgskh4elQbX3w5xKrD9RJI8CXVe/BORAL8YbBeJa2WFzavFvwvjkZ2r
JXVeQjrIxlGXVDAQUMhJrj9lsCV8jNUASOoEGus1I1IonWnCWl3vNHnc3LO9LI1c
OpXvD9WJ4HuqLUSdKU+RBdEPwZg1+oSe30WRQvfXTEgKKb8Kp4iCJsEsajpqS+vz
UEAUsTwPMGXR9gjgMEJKlVWiqupcVeXBVHQuG/XxPJ7TCwcUk/hSZoumzDrD4k3R
LU22+qbQEnbUOEgVCwF9f71c5A5Pgsnd6J+z9Tdt0ExS1MuppU2y/40+3tzVSMEz
itGuB7qF9b459GcbkvYUydumHNCNJwWMtQ2i70zVU8GIwEdLQ0t9IW4R44mCorEK
jA/lmbSDke+ausJgaPelbjmPLSWgawnQdmrAP1FkCh310GN9REZK+A4Z+yJ3/vrB
eAKCcKFIkSVxtBFQ8hwJuu6nLcIfVoqHhcdqlezfBmMN13Y4AY4z9UaDgHXe4iAf
kr+q04GqpHAP3itCAfNdxBvztuSFTanidfpIciku8zjq5mSTt+cTUJ4zHIA/H3TX
oRRUbjZno9kM73lLRCgCWulB906RB3uEH3o310bTCUzq5ucoYpn4Yqyk3ZcZvu8T
eTF1AFwaSM7xcJxgMYm2vj+yAvKwLq7p/Uc28TpHv235rctjjewZTT3chYLv/SAH
wWB1eqOPOX/7tOU3gq7YG/qK1lCspOscc7N/pkmy/a5esMaMlh0pNtdL8//gYcCZ
JOB774jacamn+N2K9X2NqPZCJ53z179yWT/4BeLUnM9xOkovOpeoDxR0i7ggQO4C
ufEBhHpSWPc2jKK4qbyCiXjIV9PaMJNP+xrHAEK1Q5YAfxvuNfA/9o2kLjF1tNv8
QfhJS3+XnPyMbPk4dRhEZY+XRPiUdoz3liEUPjUGH9vtzDBN4DZSIC+rPHp7YI8C
ASCs822FreRTIBzlxR6B7x7VtiT589jHKreRbKkmuxnuREokTmjcG3J/gSUqLkMV
J3D6DdEoMsBqC3njBgMjAAprNTOfBeLIrkIJSyuMMyM6s4iZpqIsVZLRJcaYytTB
ZMgpA/cG+gEUYaoYSwZYTdfQzA3fb+xekvQWOfbzajtDBUQXvrKYe8gI+LU2L7mF
ZJLuA9xVXI4PFWBWfVDUmHE2OWVCr52FiEImzn5A1OrthMKOsrAqjXAtG2/bWxxW
BbsDQBqxFMm/MLvCVeIBQFgb3j0u2u9tiJ1HiSJeo5QtuGh8rK+ZH5LcGvWwx7Yo
sFSaDd8wWW35G5kwWoMb3VDVT86anVAuJR10iJkzKV9xHpilUAhjpPP2M0Z1PSlB
GVr3uWcsVKd7PJeOjT2ljD2y6oQ8WsdMuPDwHqohwhUfQ+dn2o+LjhaBBX/b+85r
7kUYoP7X1B24q5j/KxuNIvbqdFYh6kP0jICCtBfvnhLVuAT8E4FzS0qlQfpzVL5p
OIrGzA/bqm76bA7LXCxI3rkCSVDss8QAE2qVB6dB7NmtPg7o2ZVPL5YdFBCwh9E7
//lC1bUwOnkqJRLpXsFMHl2A08hUXO+eLFfJ8vpRcHh/GFjC7bkYmv437P6Wiy0q
Ff1UMhATsHs4Kf0T/sUQGpJpYYuJPLSuJCx++7sbp8V8AoG1hJsHrvnMTcNnfsxK
oG+wz8ssC9IWWn6uH3OIcSsnJHMQDsr4lfrLUcQXf2VC748wbj6VeY8ORWxGsy7t
R6TqkrB9Q6PcxPNawDPA9w6AEr7KkY08sywhChcVjzfgaSkgctyfMKcR3m5eSCWI
NCMHDFoc87Zg4xg/doWANOHUw+VE4yo6uCOFzQWiIr5Ec2gul9tP7TyNk2Yfv1VA
xN2FhXckSITG94BQLoVvdgU92JoMVgmAqJsZZ4rBkoAxgh8hThhhJOSCcnzOERO8
eEBXmdUHxI5dOUPzeH5NVrQB+AgAoHGegdmB6PFN6n/D+8xMQbkhw57W16DOgkoB
SGi4w6/3mQhdhB9Dpbo8yodZxkqiCBYPDYaQlxKmntm0v3z07CF3IdSpcBpzA7d+
oCJ9b/C3Isgo2RGtPIhwmAp3zU865SCqRKGSGSBhNLjBiIklJsaoPnIXIAV3MHsW
Uj2eQ7KNsp735trvMBpQhyTFXF8LmUivNnpDKJR3CjlzKHyAwhotdc8fzcukaIRa
daUQDNo1nYRo8+xDEU0kSL/oss1Acw2m1Mo9qBOWeY94sh8tNVa+C5/roOp9eaH/
37CjEuJhI4Kkm6SpIxOp4xggSPTKC6qWRgoBxYXevghaPlCEuJ89uUAguEF7We6f
xexsmbYvAQJfpAHgyLoSAoi20pQtHDe6xyUMoDyQmN/D30rquiOwfVfxYZtdk5in
ZSHSvyP8HMd3YG+e+nhGBjDk18pWHmhPfQrUdVY1ZYllKb26ihb+4OkH4k9SxBP7
hhEEvqIa2Sch4t/mv7NZlmm4aMNk2Mk9D05kzLtLcJGRTjglbQELtgEZ9Hn66W6r
wlTvr0rqE6kqhMhIPjyCvG3DfH8crnaJiYDknCvzCBQ3RrbhXOONt1M8WzIlcZWS
VBz5RNnWB8HACc5GThgjiP1Yw9l9efuOdPU7lZmfoTH61R3jmu3t0UTcquIMV3Kw
U9oL+tQNmHfK5IxUmJKWKCRSEspswAO60pQoIM32FFejm/N6FPjO714GmJsB1+8J
su1p3HkLYTk3LTHshc2hhuYNWrCX+9aiDMoVdw7y8j9V1wu9JQ12GQfISTDvx3ds
950i12M7Oe7PuC8q6r2ZW0ZmU+RtoLTsgPAXZSvbl5wqcjlZ+xH6yCIQKLvDwUe7
q8rv5cRjZEwCxEl6lXTxnT5Qltfj9/OOZx5lSpyRfoYVQQyuORxiQCNCWbNo+OzO
tl7kSoGTU/lTCqkEuA0EDAXt6RJ2FwmYtZcQAEFJf+22khUJH8Ba/BocyrjZR7N0
8yPoTsyIlhKPfBvyPDUH/ioDFr6ChGohZ9Z5H4AsXxqHUCYy2LVi95mk6+xzMFoo
nT1z/zkEa8Xqx0XxJPp8V907oMIycYDCeWMUETNPYYVJFpOeYbKBgSbSXsqf8ABJ
VURCxDlDkMu6lzR5gTfGWxtfpLFDEfoA8CuYIfAyLlTuVjnfDHD76GHwm6+JHOEb
3r+HqV4BKfzM7uyFbMnCekOCV/Sf3vso5vCeUwQerNoMe/JvntdsHTKFmoO2CUOV
dK0F5ntLWnnBaLXpDuivl9sgzPnhD+YmqlPF7BBFkbMUT6hcMglwyslex5oRO/fa
K6XL2Xc87+rVnSY61NnQTjtxJpUd0znnbTELxrxajQcPO4e5x8pOayrt0jaz5k52
nH9GOSJ4/ifRuX8178myMz+LYjMMCxbrsIAF8I6S1l5l4jVkGacdm0ybgZlA8KbT
I1FO1p1qZTf3tBN4q3rUEarZRZxd9b/Sg79ycvBOTc8hQwr80SlQf4Q5purcVIn/
TVvAnHOoXqDv1fQaduDWxpCAHjmUbbL2MOlTKJDCzMOON2XUYKoxNs88iLVgkP4p
hSDdfiJAckqZBsbrDQ+1CQMS22aTtpDYZbKOztb1S+2vtCCnosQ2NT4oXkg0c0Vn
yGb8ebHTWc6y1qoOpFFeyDnqxPoCdhcJEtyWPf2beCnz/XBMHOMps6BAJAUj4NkD
V/UAov3Ftzts9ZkqrFCCkivYsBSZH+0zJHn+T8CXtbG7+u136qARfNOmiIa+FiDu
og0ePiX0S4iiX9/Zi5rkJD/FMJdK8f4twfap2813eIqt+n2koCppkB+3dAsKg8+d
GEXVfnvR+y0FQ9C7JXSaj8kymsv1aEIXN5Xo9NPY773tbbN2Gjs4pBG1itc7QjyR
7ND+CPR8zVo3O4dULuZ2YZ5h8YClw7RJgXdtHRrOGx5O7an4hM96a2PFWy1Ppj9M
6HJXJb7H/gkD3loSJC4T2rrwbDid57TvqHI1hsmdglK5gcI8/NJ1zmWcFFrkXdVZ
mI5ELt8MhXhFDnF4kNo7X2jO+0H0NN8SGv4No70JHzOF8j0ADoKFUP5JZ/ONOoSb
NaFWfdxHfnJ3AwD4miVa1IpYVbahIQr7Myz1PHbH316TqT88KNeKSW4wItf+2Tnf
04Gr+hs9i7KuRNsSmn1MsfrPCQ4W3D2lOQqQNKZ66jFIDZRs0OncqUVkX9PiVdbH
5B6AGxPv6KMcdRwK2a8E2fl0Gu4XsgX3jCaX1tPm2HtlUMcTjc3g2G0cZeiZNgDW
3NQBuwzMi6W77Il0EYb9qCv+SUoa34VkD+kr0nCgrD8awdwZKDk9JIaUK4AcSCGn
rhWubjsR8eTmkuIv6CjVZzOLyUHGkr4TdmPDqEX7DJE9uKxjJSBiszS6Eicu0Rzk
ytAzKGWrMjSJ8rhEYBW8zLbUad2KIoSfOZ65xjGWABXxUHh8jo3nmo3mPvfEnU7t
ZGpCV4C5odmNagwAjjNhbdS2wcdXhALielJ8tpbAi8e9rgdko6PM/IyLRdCuYLQC
ae7GWbBrz3WRK98EYarNgTMaQ2nEpD5R+OnfsZxW8k2StFp6nThro5DBUqNprL+Y
9SxkYpgS78eYedsxRIa5b+KxuJdWfC0kJakMHtEwKRE5dAWoaX4jIcsKxQ9fzjzb
wNMpITBtPqnm/iKhZsDtkCDChpphhWiu+OblIMrag/sWLIQfazCZIEHK6WslUIAd
S7TD/R2WjT9WuOfArzX+22q8VMdz2rkAWqD8gZ5HfXgxPzenRSfRYxmZi5ioYeae
EJX6z5nP9n2/7w+Dj9z9SCsgP3qX9N0f+mS9qmyELLeiSr6C/0jT34Znc2q1Yxsi
NT8DiufWupbRJzm4512MfNZyxiWzJl5VNCQQz732dl2mQwubkF9dz8KogOj3HRqn
SVicOw1L8FK4x/tIjJBKlK5IhAfFNVCPFvD5valT9SGQiJHcFtCxwzECKqO/JKjW
9YqyH6gbYsgQioEGtT9wzBSeMhNilSgXY1PToB1MsLaQIUAXEKXN7jVnuaLHs7PD
4PGn43fL85TowgMO9B7iDDtwL56UFCkMf3QATqDyiTP8SAReNJwqTUHQj+30KHwm
fTo6vrYh8zpagaN74pkFemj/DPBFZ23/CREB1EYKKQix3EWKX3JawykvRkPIgJ2R
Lg4ANAlOj17bVHmyNsw+u4q/dUNg6nnofwMwKm+gbOJWtspvsgW4ZmwlMNPq8a0M
toz9KqKRXSCKrVWk2JPGefeXlkbLJI1Ogms4NbNccChsjf+mDuWOMjKtmF1mR898
I/mtbMr6KAglKUeT5ZZ3m3EZRBKIjCLcz7URVaQ2f2Sijk4ZgeOgN8xmJuLUjgiV
jQYXOem5nT3NfdUTeT7iMg9MNK8OAPVpc+c6NPW0/Svsbi+vDtzi9p44EdTYcIM2
+NS69bvEUg9ZDuRNq5vAjX0nMsRwCEXHoc+f0qR1hewHrzurt2p9A6fu0qc4TMFR
KHm/RTdT/v+P2K16r3edFjGUVcJ1oqzZlkMijBQc9N23HK2bJ/DKTE13hYEDClUW
9rrN1yNS+70qqJDIUHwxTosl4Y9vG11X42j1EhjimhXSC16DOVwqVi2NRlIKQQHN
KEwJyUjirpFJ7eV7Nym9a0frokAO6ygBUAipbJOqizCVyG48rDA7ECZfsaQYt3Kc
0H+rYA3sM0StaaxeZzUNV/6shjT2QVyDhw1bB0dtCt9uBUJTbz6zeiN5SrXeBzRC
4D/JE42Dqr8fznHrwW3VIfk5P99VYL9G7+TNTJ4HB5cUQO7La4VjkGjLQPF0I10e
UAQG2gKcuFAxv4O0HHqNlMnTC/Tpa8XLuNdH56L5odjbTtGEMJvltArtJ0t5GgH0
1e43rLadM8Fvagwt1HkTS62Z85sQq+mITR7jhP8XUBuOm3r/loS4eylPqpC28b0e
FmcuV/d8z3Z83Z3/UAYXDvxaeeqrJtQN29bVnNa2xgoQfBZETa1nQ5XrAelpGb4S
LBqLzCTeWTChkwdxXLaZoENCqyxxTdYDktxSJBy8EbpiO2f3Udidbxu52YGKsjb5
nOrLpfcgN8uDDz6+eR8GY0MVtdPEPA6gBBxZVmalr9+x+ywdt3BadWl7Tj/5hSkO
RByfvANEmeQxzP8lS2NjNBfisnoY9ljM47k7H3bz3k5f6o5/CvE7wz5o+u9/5tsu
POrR5a1l65IUXJk3pwJakFCiZiqj65QLG3GeWuIdJWvJspExU/wgdOsU3X//GUG/
0iahXlZ6BH821vEJyWCP0ZL4RkYJM60lk3v4zd4+U125PEvEdymmaMr6MTsQgsNJ
KU3zwoSz4LEHNm2HOAVLT9ysH1D9YkbH7WxH77FfSE5ybKFeEvemegdK8mEYtnWQ
3LBZhCoLSfoTEWHgF4oOw0f0AKwD5kNcfOrqs9iJKfVa7EzF0RTCUIODuriN3W71
VD+LdUEzcgF6ObhTypT9iW2ayeDkKKhDzoxYJ6GDK+e5la4H0CYJJramhFkK90hO
sJdCl0oD/H44tmeMdLZbLj3h2EJsmA+4N4G+U901HP+TQJSGwb5Z1eMQTwLAH0UM
pjYjF+mi8B36GjtdhP7y93C4aFaqaXvpMtgqCCxAfGrHNOc4/ExFMtyhAJ85GGCV
uOcpOq1VU5KTdRT5gyCYdlL/+3QtMKgxXuKS7rN2ZZOgUhnaKqAOcVz29RQz8RbD
oJZKv7bBapR0BHmBQtu+BLADHGKdUzv6tA0WXO4+JyaywhDFi5wDYbUVk+5gJspg
I2T7DKHmz37FkvEXBHu6B+prBAbea4OfJ8HgZ7xf4ImSbpQrJjbEfbt4GEUNANQK
uGcIm61Y+uSJV1kIH+6V430cpOFJk3w3Q1LLyRl8n743lzAJWjIs1NIaNuvuhl1+
8QuxJ35i+8cBPu7t1eSJC+eWLCz6iKE6T/C1vVzy/rpvj0sGtjWBflrQ3rIzZzYc
VxOlcASxbuS/D+MWx4+E6zlUNKoXnnD+FIeAoIP/Kih1wbV4V+59jOT+AbSaRj7v
L311bUGsPtwHbUoigvfeuAWAO5IEDnnVPizpOS7V8ulgEpf44p1INAU2lifslJE/
kiOQjTxN8xDWDAIJ2U5CR+Je6rAgvniOba9Fg1U/jfWyGRt9p8VPt1MfJnYDHuoL
YnqeazVG24R492zg1K+eGfOtjRIvRqWclOmPRpZtxocDRathrmR1i0I7znOkVp8O
HibG00ynCqxYyJ6Te3lSq2gr3bZA2Fxu86Z3dmhkog3kg0a+axdGLSwSFWDM5Ill
f9VzcjlLjHhgLyKOhXD8Z2DFG0l1AmVlk5cMflFcXxRcjbX8DEgezHO+thh7ghNK
sZsO0UZIFeqBaJ9KwEHiAHVEYqwskg17WEe2PUAU+scD3Iub0thjY5diSiSRXTow
QE1kXFSEx6qJ6XkFELpMBAlO6xczmP8sYmooXxCb3dz2l63l1jKq/Zm32cMtORdk
mNEmi8XPsPbFI9bBrYfqB0xe5mRSHJ8xesDJ0NDORv4snBR1XfCR8WrrxxkGZJxT
AcgyCyPd0UMMFSTkvRozDe8H8bl7ufnN0NcNIppcNjKeAW3Dg/Vj/VI9FQBiAgs0
JNy1oeulz0DOGUn6qGAYtNuQo+lhdTdjwSWehKbMr1Jy33kXB0vM9fmhBwul0AqF
P7CfuN7WZKXims8tK6Xip2Cx0G13jWnhUv48rL5xocEDc/bNX9zAxJQhgTWkdu0O
3dDd+aYdc/awJRmyX5RJR6of80xq/meQRJ6btE/VpZQpYWTtSNaZmvSzphljS/dv
cIdHHXodDpWWCfVflwgxGjJwN+HUb5/l5YgCa1d5G3xFt1XOzr6Q2u4Tw/biywwI
v/Rd9MZW3/QRX3JnfHZNapt+8RVl0kJ0/kfNXmUXv4sDfuNKv32SRDZ7YTq/beKT
iFiIf7UdRvKMabEmgR1yFwZDnAxW8UvsIeV0C0LZUQWeExz9/SJJTbq6NNJwPl/3
yELPLnIAGSAExX2wmeFbRSu9b9wSlB7cPTEMoDDMVRxq8WTPcz/m/wPlW4c3I22X
69x0b5NtGFeTahjeUJluoPTL4D7WpT7XD95PMcNgnNluzTCN0NJaY4LY7bhLCvyj
xPpNcy56GQXl89RzV02dENrXEjT8XkPK/h/pgmPLk9TS8+U/8HANe4GR/O02ZhR7
XOtPVH6lbLxP6ySL6ztGLBGCkBFiDCAXott2YkZmaC+zCytaDZEB009sVKWH2dQb
eoRSZmUAQdHrRTs04sg1fzMoqesmr+xkdwucFvVKL2bhDuyRTN+BdmKEgcDot53K
nBZYUHg6plSESH0I4uoKlTbfbOzNq9YwoamlqBjhDuVKHJNa65nUnpHE340kfwF+
5b+6rwG1AqjwjucxNOESkHx6+oLYtLneSf1ZFT4Pp6O59T2txHtk9jZ/2EhVRBwp
xusDqN352BmEzAYKWdYA/AuXpxi7wDs0S8gyq+L1DFpCEi1PPRN+V3iEGIRArr/U
Ab7Lpm4D/wRl7pbdx1dx+AHMCZj5OqzO67QTI6JESQFAKfmYdHNAwoh0SWXT9+tb
oML2fTKoC6VzzKeyGYTqGbuAbNCjWc8jJlopWNOj3Cbn1tXoxrWIcknSk8PrYVIE
KqVfuaqTR9ya2xfbxH2uJMTiMcZU2irzV68TI6RezFujjG4qizV7hUcTnnGIIE6K
ZfOFUf31qIs5T7rvmBfn58+NUWaZJXh5Udz+VXa2Wf3xrovRSQO4NqfTVDcvBOpd
1dPZqmIhAl3d2nvdnY7jSMBrGS9uDvDj34BfhNN2SY6uKPlaRzvu8Tt8GmLYysco
BsokWmwaSYsnl6I2vobVRW7QtGet3nW0KI7FWIO0xsqgJCN5gk1SaHlx5TecrpiN
rYekCUdU1tj9m7+VoXw5dycpj1eOYKiTybJJhcsB5hVB+95n3SCYaAXxeAF5w4gI
IS//Z5uPsKvFlrwdvcYwbe+UlPKTXWh7EEOEC9n/TgA4jVA1F52+fEref0cgJq71
AgYYR6XkNeUempmwFVPqPdmHMlUxK3+dzI6QxYqzvzgXSrJcim3Ydg0XD7N0CtXR
rTcWbtcddOJ69p4p4+T/H5uvLhAlcvD+gltPM6eApwG4AOALaefX/jLk7y7lBiiT
8Rr8W5FKioggT1mNh39ZkDAjE8etbd1i1gCFHed+zjAg6h3PB4RK7WEwNDXgLNA7
3OqcXYQ17kDBcEkDDkma7MhRC1O0O+UTBcNLRIcphhKoN5Do3tQGXIxV7k/SkYVm
1awD0s2A+rFRfLiWXlcH3Z9EzUY+O6M4xE5Zci6vSXJHI9RvL2ROxZ717W4NKaHY
dp0yr/svSH79GnQHKtkxbp7olWn0WFivGsDWpC/v/GCP2FcB3h028A1+u/gBp6/f
/gIbhUP0hw43z9gXsEm8rHq/ceyW2qY0n4DOYKPLhbQJvdWnD8yvOJALm04Pr3Qa
cptmNmCvlqzaXsEYs23TKDutNkvuQaL9oRhjA9WUXTDGd9mdIXu3WQmRTfypYgS8
Pk1h4x586aAawJYTPAcxysitpw2X3YX5b6F3VHEM1Jeqa80DY+0OYffYIEAxHZuJ
8Ym6fSTcC0JJvgAIPlBDoZm6NIjxXDhvphUMfD6m3zTVqjkaMVDX3Yd8M5cIsln1
9wpbmy5bs8XiEN1IXEpBP4KwG1Ryhx1l9btMr/EJJCd9m7zS8ITeXv/hVRG5XMQR
BSfuSXAc5MzxxUG7YlO7bZahXpc2A0TYggJC3Pvilp9wqECIBYHHlpOp/EYItNO5
r4Kx4wJo3jLp6g6Reo17KtlD4TM5YI8ajQy7jSp1PYmKlZsrheoV7qX9ItGhXmRn
YgeQ6AVd7419oZQ86S3TqYMAGylxlX6fHbA2eCStDeCefZF25q2ettmPRg38oIxS
TjgP/fv+zyzLfM48EdGTzUNBiHjKGQWsfHXH7P/P8C/mEC/gSmecMoBAll/77vzF
r3VZ8Z8D5ue6HcBc9RUSIHD6kae+Kk1YR8bmh1p2/yEgY9JtWeEVR2k3r/soSa05
IrNRRhewnZGtEfXveDvWf/90ByYEY+fjNK0ZfMhzey5SlGDqdUbaFE3NGsHHSAtz
5jlAyoisK1oTvF4X10vP///EBTNwb7yhDDzIx1nWaNEjvGID9CeX9fFF1MmddyFs
TG1ShZ9mr+VqRhrngPcN2dA3X/+7daeO5PxdkLry8woqgOIqwUm6Q4F8UDAHJlP2
clR3pvrDw9iv8Uns9geakcYpreq+ams2QOulMhOcDFmX6VBNaQJl54zhA0lM2MVJ
5n1D4R991nQXs0+zhrVF6kyC6V+1sP5RiGHkrukTXTywASBnA/rePppAoE0ei3bE
IoS88q+QyXacSdDzSdKTNHHULTwXAOnzeqhJTpiWY0rYVgHy2x3E21Xw7jeX+AoG
sj0M/iqtbcFp+rUm6Td+v3gSO1KSoCTo/8BCTO8uNaHFJij6bfyGVfBC3FK4gScO
TzS8cVCwv0FxHJ/+0A1ItIOYXEqGnfqOlgJ3eulZ7Czi/wMrC++K+bgFslgtbB5r
WsQ4X4v+iqtHHc3NnJclA/U18cs0/18quJBiUchjMDExRpuMh5wXt1yn6e7cKmLA
Db/A5cyXkGFUmb1pi8gup9Rb893gb4jxKABbFd1vsT57z3avquLV4/CY8uTdV+2W
+vCUajzEQMRmuNt1Nnv22l9kEChR1VvsCIogivoX32yysOd+70ape6FG66O4/uAn
LpMruijy1tcZ+N0/s91yoFaqxuEEM/1G0Tmc8Wl3lHI2mPWg5Msw8FT3rCQNpwXE
0EMXzGu7j6RFUbVcll29smFVMRiEcXCbG4M+/nUsR6rITBePwFyDHdqUzaJ9Lj8B
wvDVNDRw6zop4ayV9L9eFH+vCsiCo8+1bo9kO+v16nIh3YzJZSUMSrWDmE0KfCqI
boDQft0ZQH5NXe73vYh3fRZr/lksZ0WhMP7bnD1M0XpTrLLsoZ6q5Aqh9Vkfd363
K7oXjRBfTq2RWlmO3gGFzUDk0s2Mj+mnW70nMKQ/P18mT3S+tep4BZV02R7eddkb
Cw2EWljB2JcvXgAiJH/1YsDkUuEWOtaE+OXBEaMq2bUqwIb1Es1TVKrB9jJdStdo
J5hZXDc0iupmHNeW7MDNIS3C1PzL2yigDi/b+BDugINHLEhk37kfbRLlgaKShy0f
U5Z+nrDAGiFF9/XFpL8SwNPyuBor8d5RMgFHnxzwH9ExtZEMPRJjhJHojO7mnyV8
vbXZXwluFOb6zRV8p9lYHWnYA2SwfEAD837PkgqljbJRGIYGEbkfvxHDJrIz036r
TP4a0ERImARVza2yJ853w+JhHvLfgPe19m+1WkuQKiflbMCSG/cL6VBCCMmaNs/b
i3DimggBSv5vj52cZZX7LJCtEH1m5QMs7sz00dwW+6s3Tl+dG9oc9mpuMI8Skj6p
ys0bH5scm4KizA/UX0MLETEBd0mC9dAhYsiqUlq34kGFpItxl+KWX8ws/fj4+mo6
z9UsAxOYGkf35XjS1eR2fFDqVD6qVXbO7BgQIwkFF5SMcwhBJVVKTee40dbocPr8
QIns7cPScKovGZryAAM+DDRG9XpLGC0qzRJpfRIn3c7BTzs6W8Uda+tIL8zzOlUy
rZe3+utNK1LqH/kSUKZJwKx8XUGGKE06oKqO2l8pjsQqgad+yBrZTuRlz3JIALqa
zi6ZrPlGxMtX+fbysTHmxTkaN1hVVOwKADgWbuFeL3cJ5zNvKKYzql0iGPiOHO+a
CxgySlC2ey1CPsFVslafAzmYMaoXXKX0GbEpW4E/5/1+zZvWvkpa7rGc0SGDsJbC
eNMpk5Nm5xs0wBuJGc7N1p8gHPIBf1om+GR8EgHOG1e+f0X4VUzGqF0AxnGWBzvu
jDTMdJLyQ4ImsduowlvmcHW/fPxDgOG0OS3qL8b56FP/jwjANK2QFYdKwyws5INw
Y1Twhqp8bT1II6+Iull85M8DFazIIbQFyudydl2MJa9W849NGbhv/LZ4oNyZqdQ0
fGu/wV8THshzpnrvuOXeAl+3yki/3E6tb0koy1LRbs0HcLhfqNarXe6cg+su2LUh
7dZ50oQkJpJ8hwJaCXuLqIr2rzUP518u4RHOKZTi2vJT1sysTRxu0PgXMw+LOZlg
wN/6xhRbdZRRrzBMtT/C3cJau0aLbhdC5tUoCzrNCXPgpAJEOZt1h6cqBs1nc07m
qxUSeIMMcF8t8XPpYECg9sCKaBMdyotfUfJzI71yNCsQ+wfpoijnMHMw7v9dJvdx
0uWHl4xxz6PI9pKsOWD0rDvPUfXv9KWniKOUh4mtGrGmkqOe2H4DJJTBb39aohk2
5oZb/8HPcoTttcoO7ztnG/X6OPYcEotOKM1f8/xzlKEHZlBrOZToUZARlPCMlyna
WpSws66HspjvEO+oN7JwYoA1T+8KI/YMNgN3fkgwn+8VwTUkDCDDDALAjjRCoYGC
0w2+xGzXARnsgrhcs6dtTOFwUEAAp7MWCo6FCnp6rqYmcKP9rvdPs4GlBmHlchuM
aWbb6NnDOAZNlfgyo8OQyY8P60NaCBucyFhcYK9gG8xlXhm1MYXOI0KRMy8+7YRA
MfskdxexWtMgJllzB6kInB3i6NtNm55hVxtJPo3bcKva5fl5CrMREHkjZpOg2y9A
mJX+Rgv97WoYkCixa0BBlVfABg5c08dLY7L2eulRSXQIwvi+b3g3mMMrGgKNK6Gk
6CDQCb6k0QEF//Z1n+81bf5IJpCSp7ZPoDr3dY9s7dpG/1C0hSRzyCeEmxpc2crX
tD0rJisa6ukHyK3IXTuPY7mje8rF8dU9qqspTcbeGrKecfB9gi/2juIZFwoAAYnf
CeZI3+3FZ+pH9FmE8GRH+bQSMweWpX79KqEXDeGMA+2BsbO9I2h+tehc2jwLxkw1
nP48Y1QMyi4CelF8GLJte83uiaMP/xyRQnrBCpZEHLva/sbKQM1nVejUq3EngSfJ
rfqCHY3MEzpnhAViR01iNZlJ0jAJRdNW48ium8xMFdB/j+NpqfOdtA9/HuZCY+ge
35KAv3EdezSBm6i64M8sj95Xxg9zILS/ZkJ0s3jO4HCJTtzuxgRNRkdVLIysM1Vr
RSJGa2iFPkcA9kVNgkuQ1lRK5bWXt9GInmQ0KlQgf8Nh2JHgIFfpCM6l4eJ9DUkt
LzFcrT7UApkTkBi/0jjdxqrIz93FLxFvFYq+nZZ7gH44dhqo0L2JqgdbdpMUd8CK
KOEbXek4cZvv7RUCvrsEZ9grkxNaokg5BRLZKYm/2w0HrDVSGCeCCHFLzNe5+XNN
lEohY05rdt8Q+I/N4XaaTfAWl9wkLc6DBlWlHXba3bAp49MB+aOiMgN/JB7+Enok
r4dKq9HFh+1SluU0MZsI3mtAyTTbuLVo6dYbrbXvB81tbdwrTtX3uABz9jUDiu9v
Q8WPyRob+WssaDPDIQIEw1DldhAZZga3qw8sP35FHq/mUTxoJ1BUbieax0DGeYiK
mzAkOrQufHtRwiIVD1kOozFlTbQh0ZqlaeVbIXAnCcFf78ayWy7PyiXeooNxy/05
zL7u2f2xuubl6tYLBGwFjIBO+RmlnMzgbupmCClX69WblYnfLXUDXzm2/FXk8v8A
kcSxKfSMv69bUaNyIlcGK5ja9lhxqi/XpbUEI6twWof6Owq/mwahIsK/FNXv+d8B
MXsdctfFEl2DAIlta1iCEfi6REko5JNY8Y+PDnEBzS7MIoBmDnVNLdmKznpgSAuM
4WJIRrYdCnv/yS5q32+NyEZnEPAd2HAxnFawJdnqCgSxUbyggZKAl+saabeJzk2h
NmJsX2REy0pvRdVkuoS8O7HVNc8W/S+enfjZBw3dfLAkCTAIWvj2vbm5AgujMUf9
+ZDzTSLuhS6+swKt+E//i/kFONslrkhl9Mkbo3vgX4UG625Rqp2RmPjfOFUp+bem
P77zeGjBMY7rbi73/SNlcQpvQrTEBLfDDIfx+6KxuaNorzd+ghfJo6OA8ZrdpF2H
NvxxK/lrgzzKEUvv6K6z4RklEXpSzjaJg75mKmUeNPFW8CFU6sazSjcdxR9Eqwc7
ZdgNxfwUjcrLt7GfQxSf58U3OfIKUiDRYg3ECzIvEvASrifEMAsprRqcYw13cl3W
GhG+Bw4k2XlcdFGGgYiHVsjApZsG+kfbSeuWxvb5ys8VK/Vn/J7sMuFS3EIEVucc
7yCIeUbrkTEjd4BS5ucFUTrO+cqge2OjdnubvaB6WBU6M+AcgMsIyGDIsEGKh0c/
GpoRhMTv/HkGxTEAImA/8K3WuAbvHujK06ooP9IdRWcOe4vt5ngTFXXteYX+BTW5
JIqsLD36QgHV7DDFenoFNt0+/nte1rFlM2mjLJia+oKKAjWbDnCxsmTFqhzgODmA
iWwpWNK5yEhwl3MyDTZcg0qmbFkkvIRbXOQ/3c0hJKBVmi9uATrJxUbpDWCBLa5X
PoJ80M5mFC3r6WUNNasi4CWbJ/Oc8mbn3BU5arOGMrEWsh1VaFRJo+L40CDuSRS9
Tg53uLR3wHSzlPSa7xmdXlDyFGywP0I06Unhc3l2drDIhJ5GWnvHqBr9QlFEKP7a
iqI1L//bQjIZyidXjsrNBS9oMxGnpWhPlE/aJvS4a+ptY7pt1Yl9x7NTABZ2eGqS
1VvLYW/PMpqx+gIgZ4orWhS0RFeAvzRxlzwkruXlzYVDYFC/T2nGeIhvQuQEcuu6
3uo5C3F86f+7D5c2y+N3BEcbj0ZK/LAgonKCDBsTMhHlhQhitOURtXUAFOU72TP7
Xwz5bDiOTvk+fGM0cd5jfzHZYu8Tz32Y4vkYuNndtxs876E0LQ9AT8v4XT8hYz+d
ymYzrLWIrMK11DEpterb7BJq1S/+ox9KbrcXv4X39pvRlZpIZIe6RfhGR43y3Vuh
udR/i0jBSdU7F0xijCo3ZR6DB1JyK21rvCjbhvWEw8X1rmKO9rIkWulI4WBBRi+2
oMd82baLmSEiKzeVlhJdEbBCl3kDUIZwLKWvRIF/I52NHSysQRCsEmt7lIdupCaT
NXplf6ilKuNM2CRP7zHRwUye5b3Suc6uKPiJ7bGTxMC9h6eaehKmvf7igwp6cIIt
cQcvag+QnunYszwT9Bmz+hR4T2t2yg7w3hZgH49KpfWjruZlZpukS09ypM1P7Sxo
nv8k7m84FV1GN3f+5l2NV0TkpQmKwPnunOT4RjEz487y8ZQjLw+dayfUO2Gu2vOj
wPkVjMe94cjd2m/DejRifyNrdLGUtNe7WltrG768/pvn1xbcHj5AcE0qL6QPF1ji
u2hiP0qFlWcrxIN7kj1OyEcjewgeVELQ8zvG36jCyiHeJtCOUWz3FjUEMY3vtA4Z
K19LtVCqccV7Ews8UtRi17F+zJwnb/RsIjq9PP73YxUW+95MJHwAklIOxpRn2BlV
OxkFfNUtheZDFyfccIrUbZHeA7SwcBBQ0/3uiHr/EGcyinwdQM2kCLL/IsXAeYgr
X1S/LqhMMuHXD/6oTq7SxSgEZXvgVroI6WPTu5MbaqubbvMZ44J0Pzho2tKloEni
PPPGW1yehjUgy2ib2dsUFSsfQKfZKAZkmA+QlLHmbj0e6MSfDrlnTqQ/weQrve2d
l5SmySh/ESppXjvhLHDZwYsxOOsSf4AB5D3JHLSsBP+bNlK4FcKmwtqBQIig8CHb
OyibO4G3hbb+WfplyfqdXDXlGk+VQtiPykHD+Ch30r5ACysAgVScrHBYGdNb0Cfw
fHgs0AHJkKcnF/pIV3kRTTNJwcYeUJeEipQ0OVSdetftsLl/Tvv39desDBYV86Vc
7NVm3Dg8hB4bYZv9W227tnQKxtT9m3oHpkCZg9HLHzuol/VM64BKbgcF+RDnR2x8
2Xd/YumrpylQAOBqGyA2mqk1ONZS+Kjp5bWL1Qu+51JJQO0owQi8ZxvEXy2M68cr
g9sp8wVQrmU+kFxRUVGHaE786PqQxUSOxn40uoCYodU0oYObQnIeS4A/k1ArLvu+
r2KGlmt4dDNDhD2HzL9+/MXfd187vuXAX68bzv81E7wcft1v2XdYq5siPgWC4s54
Ayb2ig/o+2fz8Y3cctE8KMQ2E4KsTGPVj5jhONHDE96c/serqkiYWua0a3aYFCye
xrSE1ngWr6LuadzKxejbgLP8o31mmUCTSy7xeiH8HeD1KEHwYXSf2HDv4BE3Ln4E
ADJVyaOToiuA5MPjCSqXJjQdaYk2yTb7xQjBFGMBPCD0SRhZgExb1C68oAgay1rx
DFGMnN1ez5vTkohDL3/X/AmRoxZx/IVi7xcC7yflYvmrdKeKUMgMgckvG7uGPQXH
Gbmfn2znmdg2ofAmFkriNCSXnOv8D/qri37whNUvt/msuuRc69C1JF+aqkFjE3yT
BYV6MV2I5Al4cI8r1zS/Kk9zNsa7hnrUGrIuh351KmaiIwTri1VoPRfSuLIJCNU1
OkGtDtlHnBBBc8sMy2UobVGhbMk7AU1f0bMMnspJ5Op6O1xbiVTVPE78PIQ3Of6q
E87sfF7KimYcL5AP64X2y9LZR0gEn6b66u2Tao/W6P6/0fWYIrNbMWhmR/wGfCAm
6HkDirnrinOlBh7KjgXa3uBYuGSzPNpFc3qdyUKMbkUuX8Asltb9WsTLNJ1HpBSj
k2a1YYJ5C7uvKcNdBCNHh7OvlC7eFovXntKYyhhDGoClDtZL9A7uMuJmgBNEIDIS
9lXpa+GE/g2fds1B/VatRTzyGw9T1YpsYRlS5+7az3Y0bNriO+R6k2y1n2RQ5ddw
HTwYE/kZZD1OFoOoeLNbGBJicggqHhVKHVENe236OsKa9zM2kQD/ic5uts50kulM
ixeulfH0bsDvDhGjHjkaHnRuTFnca88jwRZ1F4Bew97VJyPmdfYG1j1g5wlBEv9b
7qeFh6lBOuEDqggxMNUkgZVZAnwW/9gCxKlXdQnOu6XSL2lt8FkAlckDFJ8FDtdh
x70Gl2qMiP1MULSWc/g6ldqd/rQ5Cp1nDsVse2a1QVSXBihjYAOjg+J5jvbwBciE
ZGUNBmzkNfhGxyexT+IjlTwcpyvEdQAOdNlM6zBoDhEf0EDgJQ1J/VRTdlTNETE+
SAAY9L8uo1Mxhkcn12kNf1s3ABoSnK2j9OOPoneXKuFrveMn+mlK4Pq+cbsvfhX5
+8HER8MeI7hslZGuiZKiBFOH7UcdToM4Dn0eUJrXmxEL7SQFMMt1HNAIlMmH8QZK
81q9NxhOtrGB50yPdRmsqJCqW5Fj3a10ptmwSX/JpqOOsOVv7+uzAu0Qrgz0ljNK
wHTa9zkVPjRyBQW5+CD7A4KnV4xcyoBxDU1XqnKqHcOXThlE7tQGOLOYtmH6digK
1MUsMHOE6sz441+EApDchHYHyBcHLshVxCM9CCddSdSOhaUfX2JGnbghqcxSzCdN
LDkG7e4DQvLy6LpnXx7Vj0KgT5vXef/WuoOyhat3ilNERsfEvkssQtuawGUXAtye
p2mY1VScPoY3prm5/UNyZmwZUj30IUA8TLCTm3LWTcvqnBTsqln7bkzqcTmymXXe
AbjGNJFuZIAA3DwN5urtch6tIb9YHNYp1b+dzohxDA/Rm0oAmS8SAqCAJft2cWGf
ZIrO9nXVb234U/Wu6mS1r1KwvxT/g2I/7rK17Pu5qCNxFmwkX7St6jz30SkjHsYc
Q40YCGazCAzNQX6Oe3xJgwmkmmm8AvKgvmTbgXE6ZIBUj5pGLKJp7bnfweOXXqFQ
Gr15gsCdhXeEdDbGgiGF35DBuxaAQyBPaKARvdHdLBx71A8LYGc2G3l9fvj00t3p
rqAl6d54q8tTU2OPZ8p2y9fPU+IGcWo6/XKL3qP/nBGDjHQqDGawYTb1D+WllGGK
E2/MnKWZnmPAB5wC41HLvZNafPSi/pbKagRgC1WiLq+6xhjFalUd8n83uAlxLqzE
aptsvV346crcOAtIc8NS7cIiM+hXnX4dE2h7uIKdpt/nkfSD1+K+zVlWFOpbfb+4
icgUTAy97NGhLCO4IqAHcU8I0FtdcTIrJZ+8eZJF20+UwcvXC0f6+eHKiZVH/Ug4
QFDiI+w3EBKj1U59Ft2flapnMsIs0Znt6afTogx1YAMmGXXEuVBozn/HgiV9FJWI
7OPkpnz844IPKs5jwZa+gJ4Mg74jEt4oK59ovQd7pFXhFYcNB9vXD+9bctRFkIcN
xLRG1TutP8P/PT3f1m5Pcm+4LC9kve4i8JRKPECH9jXl9rXG4UDf54C3tzn5bXco
ArRBAKqaAbMawjjFILX2o4JJauTJK+ISJvnfhfw9k+vTT/RLkm9UhrLU1G+Tvjic
LrJYwFLj0emljwUNoduVFIlBLOzF5+PE9rfSYOBUTuBVd/YoIAhXfgpAsU3XxGlK
kM3IG7ejuXsWsrx7UyXxkSCvyKD+MT933W/IlA6lAnQhlXkEiii7HP5MdWDGFg3h
CG2DTgx8S/NACL2Y6Mi4jGOBL8TPV02MtDmSNafs+0zHrreG5f+wDdXkfKOvVkS4
3s6G7EjXRnUj2PaZ0QmJ/rEMobnhGBc4IaOyLgxkLpcn+JagNviy+wurIMX60cyH
pFvabFTBM3TswddIyRgPAJM4N2yA5jKswWUr9NSxS6xt9OzoV0hUm/jmbn5GYnxQ
mL3yt9H8fVpRBExazaxE7Gs23n+Lmp8+GN5Xt6j6wNGPQtskmZ+aw/63wWh6hU8o
w276auWdNWcZSN1NnOoAPiPnDW/F+DL38yeesl3c/q9ug5rbsQBsar5QxOkTBSt3
cWbDzs68jqrbauM9CXZRvh/jxuxTg7m9KCi+8s/VGhYcpotX2il2vJKtSe4saE3K
E4VqdCNnn4CNqilA8UqoaddRaorfxoappVafmUfZK92tEvrlQKNP5EkpZWsrKOdm
vdz11GsCUBNxZ5oyJ+a6JTd/FGN6nUuWcOUr3x0RNIctjyq9fuR4EOvIvNs7vPbn
QuOOd8MRgx8s6UYuHlMA1uuy8iikymLSwzEbtYsQJyyWAn8A+3ECHWgU5cKt43en
T2D28XCGHzKoo8FGXrtDeAYnM7X17ZJuh5AxV2MX3K+rSVTyfCgDC395XziaVWBj
854+nOa3JGAy+dMzQYtL8QDUrOpnmodregFpJwSfDYle+Ndpu5yyvu7PIOrqog4M
2RdfPDctTuVj3ktW5luatbako2Pmaz2ndLPYONaOhOUv5QjBlkShqD95i+V8R4HD
XmN5uVRD5mDw08cPvmMX6/091TCV//vPPmPJWp+q3Rmt92KpNcBk2EcuQojwwcCT
PAwqvySjsA6vAroHsTCqcmZllIeZQYPo7QCRaA27cDwxV1gUNppAczF+xY/Zxl/8
nrJi6zaCsGihaknP5W0XGaQiYK+WtgPuhV4b2V/zawXB6xFBiuoBASDDS6HEos+a
DzeMYLc2LGi7FRDAEN92QVlJhyapkvhoNvShXQWk8zxkp2Oy15+j515HiQxbX1gM
xcy+P0o9mKHH/NHtxgFhBRVH9UZme6W62GO4gqG8OBO0odzn5KX+v6Z1Sou1btmA
IGnMtbDOvH6GfGLRYWvO1/Xgiy6bbJCOimoXTvSORqhzkEpMMpti9LfeKVUUXMr3
7OEdsKbmSSBZs/r/gh05ZOwO/suAqyCSDFJUi814Dxin6bUXayWOpc0eaXY1vceT
/GjU3txMmXbYpyAhUIQs1CMXRfWqXhUiYFhkvOpqbl+4AuN/2a94KErkpAq88m8a
EG+ON3P5DKKBRaWK75MpZ4Z6nNEP21MYPEZWn2u8uf7MV56bh2V6Ya74ZMzrfygM
9S/Fqtgt+T/EDRtKin84LmX57uMFHWEamWl9MPX0IWlOQi/Xjqlh/tHn6Azisy/7
Je8iINvgvLj7i+Vcz8zFKFCx8m2DgmVR4P1eCVLHo3TjZJBq0ADta32tov3gjrie
jf0MagwyjOIVzDPrj3OQGhZ8ldLaZuNbLiPOCA7ykg5ZPHrTa3W05V3fCBmHhEfR
BA37SPPMnxC3L5oR8ka3ZhPPrFU7GTwiPN+RhJ/U8+dJiimPPBkGMu7p/HqRmUEL
0tKMM7Ohctj7eso/lvjogMmIojwtLkFZhFlJ3p/rQ0wGLJQmdA4IXfSASMl34O3E
pcpzFxuExd9But7ESOjWOaRVJi93eBlCh47cFsj5NquHlqn2NVWjcTe7C76EIx7V
jNN5EBn1szixLxa+0FAy1l+kbxJ3n7oRkbOnxRIlKSoAU3EKztqKdXcpYEK1yvSc
q58qgSVdLa9zrsJTWQx1c4bCLKRORQsBTCEPiPDM5lXv9c9aehBCCILK1lbpr2HU
oiJ7mPjaMlxyXl5hMjcufrRI9csVXaZwVpi6l+5KZoOl8jwg5iaAxYLj/is0Bf/y
jeJZycmVLTwphgLQ14InC2slAZtitzAS91hC2JDr+WJ//WpqkRGxbSTozGhdD17z
S39CS3PdYM2FcLpQ9nOoyQa/I6W9WmokgZ7i7COhAGLpXcGQvQ/mF7BPAYsAvXyV
Wu14Fnf/oRrJ4kl+nI4DIXebwlffkY3oGiz+6miIc6FqLAcxr6aTye7F5+qH1hj7
ZFKxjhvnqhvZ5qqd4+Vpz1oYidGYE7W9HqFAE8Jf8P00PXSthclApVcJuLAYeySO
oVM+I8ks9mC1pRttNA6g6mgWpm6WipKEt3JT2TYPRw5mYo3/4eGXO/GGaJVrA8dt
DXr3okuhWYAtPkGkb/gAv6kWmR0Llci3DbxltVv+7iJgyU47vc3eIY42v0ZoY5ZO
cXbh5oTbTW+dOECH4d5BAVLDIQl5tqD6Qd3RaLDuiltKz31il8lD8wenrRVHI5/0
Rf+Yzw+m9/v6ncNEXVnYLi6hy93kwZEvwbODsS+0Yy+ax9yz5eYu89JisNvLLbwz
YRpz7k0D0if9E8XAn9+NwtXA/hPu3KpFAxvQJCXwTy4PJY5l4eit9Nb76Fxr/eXj
UR/v3S6NMJlT/ixgTa0Ht6RfQ/cqiuLft5ckfI5MQvuIU13+iOQ6enhlzoGvxtYd
3HpVSD7J19gSMU0r0ilbbUjz5a0ck8KJeX6Twh4yWM2JK2KpWbK0yY0jB6JQNbYi
dlkaYB5tLRMlVqHY+MhaskOC3KaFNAU00DdxD1nkVa6UOp9z2Bwpe57KndP2HuGy
CdEdMh+pfLZnr9EsNzIfZqso9aKLxpQJtH1qXQ4nmbUA4R1v0Sx/spuiZrgjH7vj
G+F44p7L9M4SBh6JMuhmxt/TdCnLWnDBluZNBjanyXTADrErIPa95luav0NyH6EQ
jq+sgSehwSeSdbWvV/EluX6DTHnkkE3lNOpcc2OPV+DRqED0/zk8yQrJAZoLmw9a
K3fRVpNaWAm01UAvrfWjcsQ/d0VdG0XtVESw8PWb0GvEENvGmyzk4kvO2z1F/At5
DNDoQivzlKzoEZK4mTi3jYD4dOpQCfT5inFrvEOrSX4SqPeBBkvc2LZBntuJIqx6
YC04VG5YEk/9p0GROsaiqRWbUyIzW2FmIvvXWReRjlCNuk92CyFWUh2jrLXjwF6v
D/wa+VPPjwxvNcPax/Sc51f+GsRyNxE7jXFEiuYZbLUXBjllwlFHawSXb/gCX+cC
hzQZe1wiKKnuDB6zLOLn00mpKpt7S1MYq09quaRMTbENWNHVpSJLdPPsabtXtN2V
1DYdv9iZf4l3nimLo6+PeZ5rzyb/R/WPXlrErPb5q8rmmMKdlv57CRzZSTKtTaqz
KY8Mfrdi4qQase7LvsZTqEsHR6VE5VwXoGgYX8vUzKY4Ea3uBrJTkdGrXfzinNwk
MQLVEpdMz5nssKHNES6/t2ItMwxIrhIz7lpzdDb1AMZWd5zezXN9Q1VVuZJnDL3N
7Ee4LLSpRjAlJx7x7o4F/bpRzkWxiRlQhUhhAaldeKZIK28LGjmQaEIlNUXuF0Ek
hK7hA8DmzeH4HwAV4j0A017ImP1n+DrvAZdCWr5aUNWEN38XOIhc+B/1f81ihezL
sQ0jTuT7V2oY8p+puAX8mMH7CnNHNKpU/szdhHZwHuDGDicgSalFJPzEBSVPFxX2
mDqrO6Vw5mEHZ/xiYLVJgubQAnD6zQXhrDeT6hmNIKzHzqNEvphS0KAijDhAytv9
KzlfdD66eQI+rBupzYKMAu5PFXtd29Jh865arVAgD3ucjQsnpdK9Tm2F8dhQm6/q
r3sFWH+14IBWAh3SBcFldKpQiWQpwI1yr/SnIbadtGtotGVaLyYgWzFO3dqqZOWr
1L4cKbx3yCML5Q558e/qiQiLn69PLyGUSIInGLvC5sUetu4awvu2Ly33oMsebEZB
x7KKZs+b6nT6lzWsRO7r1e3oVqBnII1/ZdxeIQ3peVx8tURDVenaAr4kEvZ7FRNA
dRTNpYkad9TBnoSjf0Kwsj2JSM9dhpAYh2OtlvFdv4Mhf7rIcSi4MnlZmeJzs8yl
NVQV4EzKN/OYhREyGopFqoyEAqGsiWRuH9GdflfQkJqSaUQeoFIiPr2Ful5AmIB1
F2NTc0Pc7vEzotIe+UMDX/OcO9yiL2IDWtmOvJk6shvLl4xBL8HdtZ8spfjnUcdB
oh4djr9v6DgATFKBe8XHTqKqH5tJaiPz6TSlODpflTr4nf+hjg7RZyrN3CKCnIsx
HJQPOGXuaPESwlpSNNEn3IXI1hw9ozQakjb5NopdWSI80kZO996zFnGfbAuqyRP4
GIE3rxgkG3MS+xPnmY9e3K9KeLWOWlqa0prUZ8G6BwTs9UxKNGsaUSsLSDdrNmak
JtCrbVUTOLRyfqtR25M7ERFCy+r/A3TWTVbfJwrdh+krPAgLco086fNoYhNTRli6
hHEPn1hKUFqce6KkLZ+PG/4ORY8IGfOpf08iCdx38TLABV8XI/1FVfNvfPhdOMB3
9jdHenOeUtrK2y4T0/H2tCOvr7ZOiyBhlg7eQj4PmtJBR7ygOiAW7uxzKNkiHz3g
Vv4ddxSmV6f5QsSqEptBSpJ6jqmEFiov/RFFKYMIR+U41drX6mAw1WR3QkbRA/JD
4tR9DyzHVDQdF1i/oOHQVe+IrsrVcQ/SjpUg2la0RgezUAOA4aQWSsh8B7/TsjFK
oNu98gTk0IOlbfh6DTs4ZEMigo+MLSsYKFbwIwZdMJuw0/u09GZHdm2SJAfvXiuF
TlMba59+1uelxGDdloKIgHnPmGohrGbTv2cz7kxbGO8gZdyWO0e14m+lXVTTXvdL
+5AnHcEEFtrjdp0zau9o25MTVjVXFziJVsm7ZSV4u7YHlOWW5SaGex9vyXVDgE35
R01VkaMCc+qaxwsC87ai7x9323yXGa7sFQicTSZrEare/z8drsAn7qgqYjSO4lWw
lTPHP3WDiw9I/yIT+A6S5DsFJMZJhzGiNwELlZU2cPe5X2Pk7nPIXEfaLQekooZJ
2NcHU1TQCTU9JNv/m4ZmPwoXcJcTIASzGQiWuOw2hKVSSQZ7xycZpMVlXgCS3sat
y2C5RBWRayXZmvFOp0+9XwhUP2Q0TMW4dvjMMdZKaLnb3cWDKbNT+qmbCPMvwxjX
uVOC71Hm6S3oFHjtdorKxzfHNe897VGjpzDHK1Gkv2GfBOIRZ9gtbn24UKAfJbUZ
Ij0Leg7ylKDv30Qhz7b4YHfZkU8LB+FUokvWFHERqw9AND2mOq2e98GfsL+4SuqY
yUjJ2gX2fqjCBrASffUqjvIZYwuj8W1wnQrgHtTw2Gm9GUijnWtriko3BIPjKUlH
5hGRhmfIZ08iJvrN7Ilc27M/OWkGVvRP1YTjuWGN6UbqEIJ3w9+DRO5wLedO6zBS
IpQJMYh9WBKAKYjxcP5fMEhCgcM16O3O47jZ2yo7SI67X/plQLJIswmcjxBrQH2y
vijfs3cUQxoVZzyDn/n/NlhuOwk+pXERDwtib/PyTDG04WHvnSRViwKjfnm9viLW
U0higigRY1vdpsQVPvIEjWwhqhTK3kiCWGkx6S1qliPmRFobD/alA4ZX6wMp9gr8
zJhjYRhR8BGbpTywO+7JcWiwCTIvM5r6KAxxxtpHG4DV6oS1pYrHT3Xmo6ERHgbp
m6RKphRRgLbzKsfSg5rTXBa2TCkhquODHs29Uyy5SVE2IC2tgxDIxZcvmuUm9aCp
j9XnwXdQFc0GYVwmpfKriATSD2owCp7Yv55f0o5gNJCOa0QlMSuiR/aLK1QT0HMT
ehUPjy+Q79Sooq/S5nm63K2tpUp94IwyqMze94RBjEX6mmwacgOI9+HXk/iI12uA
/qwKhUqL9oGM9aGn1JHDrsutt3w49thVi0t+sfYGZqDrOjehmNGpr5DpbGl1SgAI
IflLvxK3WQirkKtwwwm/ZW0kjUV3yRvZrjapMEnhdQ8MYROwZ39YlhClBSQkT8Ei
EW1DeF5eP9Tdqkf3xFHEsYFjI4WKDPbjRBNrvkmGNjBlmqZQks+LaMbFaurPWxWk
URq4ovUGhBOEkGaqcor4KXZ5f3TlBH5caEsFskwAaaZKflvYgxYekF6Chn2C/MoW
oAQcObj+e4B1CR7km6e8CiCjuLglnIFXXnLI2uHwQpqM4v76mREJFGthYgFJNTR4
ZklQpO3Tl5xoJ1myoAIgV5nvvjwu1cq/JRAMdY3bAJa7aBxW0/9XN0SDOk14H64S
fFeG5dGek5EULlscj0OMpxqYRLA+eQsvRPO6yhT/5JMQgojp4SzwGt5zsti2ZTpw
rh0TCO8UqPkAqpmcpCz6DlTw9EuFrcO9IWI3nf3/vL2mUT+wmOFc2w8EGPEyLyfD
HZaXAtw8AWv9cgulsfK0h3KEx938eoRSt5hE4+lD4AXWApa93aXdfIB8360q4dap
athMR0X+VqER8EHWg2NzAnu1iW2/OgvrW3TQ4vdRahsbbwkYp5xdhHiBYNc2DMwI
RjjWPF/Bc8rqRrxA8qIac71P6OvMm82Y3JQsBFSaVBQhjsS7H0wMtD6qjBwzUWvX
E3jdIRuGdEosDqgI6rhZ/oTbqJmmAD0PPAu0JrQDN2ADzw5lZG1MEqQuJZKKSrHK
+NrT1HWW4VG2zUdqYmzwvl+O68IfspCPdk8Czc/vn7WQupc0LhyWvhpAUd6BSpsg
0cV7OmMYkon2zSXDqw1S6dF9FlOQMenyrzFRc46weUAJr7JwlIyvudbuYSZWJrCN
xfnPCO5ShN1Mm8MFHSGfl952alz/MbVB39Gl+LymU5esOcn+8nejys2Y0tJJbOA3
PUbTLoRIUjIifxDGZCDAWKmfa6ine3AgqcYseVWw6AtmtN8r09/0gPgR23qxM3NT
E+ws7eLdX//GtVXKGIre80H2Dgmhg8tR+53+WQFTP5eCgKUZi5m10dK/A4dCD+wA
K61KqvzASVDewcNSC07wAaS+BpjYJOjQ/BR15dsSYDLLgdB5yMiyvpoaXNF6pNf5
8913CbsHbN3PM3km8NoU553kVo1k2sT+tPLPS5SXtWsYuGd019yifOwgJaNJ0YJk
P+TsA+9crdjyhZE4e8jDiPL6e4/TeYFBeJhWp9Ey5UTlTMuiwsP/Xd63igj9tWd0
7XjjLmeNrqgztcg4feaXpGHxn0rQeUZYN0XZeYCPmmcOz8Vb/1bsYOHYwGVSPmjA
JJjHywHIVVVO3Mp/wy+jMbJbzkIXPKy1eYix8O5WAwV7FgDR7KISf+oPeXhq0BoK
epFSuKoO8leRKmK0rQ6foR+x3NftyDJkfixREvOAwMLhvaIVwRDhe8cTLG4T2T18
UGkPcqh3H2O/NkinUo1t132wAqfNKZ1Ogd64js+//n20Fxwg56FzgVfx69tyzf6V
ZqHKeBV3MvxScxoaVAlRkGEaUNW5w26vAk106zFls01DChZpyYaqYMxe8cB8ANad
iyeR+tbOThX3wv2polhtqeLjmyiXaFHI9pbIQe5WsgTdC70Q1v9zno04OIVkVrht
Oa32/FirZNgum8RVAsxdfZGYcbOb3FK3tKDLYnbFcKE9OOz8YLlaju2HNK2X9yrX
b3D4gSi7pZqInZNkJS3vDePUlo7fdDruGZzTepyvdKYA/jkgHGR6yxLLRiwuXNp1
k5eZ2aZN6KZeblOKm2dnSVrUhmksKYJURItaiOzZQVXIgOlW3kcMI0KjlxNEAgwI
T/qnkQJFJFMi57ZOlatrdBgm2PQlJHobzVpe1UEbydOF7C6W3A8xppXuu+jKz5wd
ZMKhMAokqNnufKzN4piTPqgMBlW/CN0Lk/mW3N9DB79OsSbtZgS2oadQGvE3Oygc
NtiHgTnR4bVtUN7Uh3DvEOWnESRDzSuzmO3JB+EF4xNuZUmWdpjt+N/e4QfaJkbp
3Ji1Tu9koUrPEmcx07f4At43qqFx4vY2T0hopC6d6z8FMTiCMVCMP1V9t4VlXoNk
I4AVuUnXOw9c3yl9cwxeKbQRucTSdSyfPLinBqm6Mb4WxZf2siE5NIhen1k5CEpB
eNDD1MBSq8b0/towE25iwrM+dHiUpe8JOQNRtxj5OUNQB29GHcJrNEnW3xnCX1KR
IO4wNi0qQLiF6qX15HQNTzLvpe0U5PPPJ8Ap8Vz7fBZt2rFXCJDUYo0E1l8wA+KE
UBSNIBqiECjIP5KdARh1rmcIBq3hQmx0QKqZsrZe2GcOyBlaKlCsXYgmJh68dleg
FFHShS8OjXeLLNNFC2Q5ZVuOBS2coLrFCNT0KuI4eWvsP6Qs1k6QT99wSDTZh1VQ
2iBuBW7gvDdksU42sQH+0geOg8t9PQNiEw9hPXvImZrCkAXn9q5anOrTcVLZvDDY
o16w169Vj294LoYYBV2SiQnkI0H9eP2uwhQf4oEm4QK6k2FvymOy7AZKExoexSGU
GsZExP3V76Z2pCegsaF5XQ3OPUkpdKYwrQvMyb8dvtpKO5kXEIKcPxUfZgRwvd9o
dhn22TUdO05fMLtnKjfkU8pMZJYHUwiaWDLwaHeo3+ebVGMy8yfzX/GROxldmhaB
36wqjFWps17MUdnir4Q7jVrt9lq3Sfgfm05gm3CIFpRYZOI3qf4NK6iiCtf5XmiY
eTC6DH01UbBYmESF2igCBuiPkfDSxEuRh48NBgZq9LwfO3fMQRR4pfWZcPJjmFIR
LSxs3H8LnAvqIOvdhg8Yw3HuSyVhADoVrSm3UpEmJAVVhWgNvGzywTfXTIEtB2A1
rNN3hAZfzb2rR/UqtNlt0IoDfRqWUtgCE3jHuW2DVUGGC8SrvQs0nI5oOy3rPlQ5
Zg6g8RLfRGzTCEoDUXvT2zXRfa4GDwUYwLchv7Tmtqncrahm8JDixMDYIO968bQd
juLseYB0JnBK7twa7HbHSK8Vf6adbanWJV8xymFZIKAImVVcYc39dqOLrO6vEhku
szmhOMaeFzVGEk+vqLKU0n3J8j3vSuMNSfCiT8/48I2Zl1NBAZerI29LxICVIpHz
UpUvv9Ckkhh6QJIPVbfU2VSQFx/fg1wogFQT3lUyGtyLm1gzlV7ZQcJpA+HZgDIC
mkFZtN+EEa/rWTGhPsOlif7YOYQF99Yxj5ZVgyTSGFLYh+h1YzfD2YeaEmTAs6sz
/HkV/dCCClw6ZxHX614A8Dm8BHmN3oxwgCE6M31FZMrIvB6R/AslSAtxsFP4fkvj
WbvrE1Be0uZxAOJiq1gqUIzJmZEJi+Qw9osWn5baFQszpmfVJfpVveCVJ4CHe/EA
zfKWKq0MV+Vq8PzQEiez6Rj0rwKi543nJ43ePe1Xk933qLqJvxnQOha+8dDnCrMw

//pragma protect end_data_block
//pragma protect digest_block
PsmCNHWfnpbif8/9/zj8Sh7lAeQ=
//pragma protect end_digest_block
//pragma protect end_protected
