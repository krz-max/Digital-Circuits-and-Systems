//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
3ixjf+EJIg+X5498AzjY55LF2XLFkrXxRpB6fjuyELjQeMIhfvE+ssM/ckJJO0dR
DMOZAk+zDc/BKw8zzXO4LMTo0+oakljuNbWVWmTbxqPxGQL6atJDYn4/6j2bKcDf
U4yraMkyfAQXmM3SqpfItuD1cpjvisnWz48+VSbTNxHnaSx9cHJdqw==
//pragma protect end_key_block
//pragma protect digest_block
F9JAwSaWlPVtBF2cYYMrMFVzD64=
//pragma protect end_digest_block
//pragma protect data_block
f0JaoYFEjCsoc3iYVUJxJkAtJk3/R68x1QPOqUdvRPp60b8FKi7jazXTv+UkWLHK
zi949kj8u6cjZMBzzAyjOcXSq5EskUzHllJOtBmUjLgL+ncWYdfqLlzOsE/Xxcit
fbDddwuRzGiK7D+i0RBUpRa7Ww6ZdwmUSejmL/cM5tSkqvHDkW0RPTvFrx0757J7
YupeaZaNLhg14wuiaptxiZ1Ga5Z5wOgGFgD55G+zJgCK/Meo9JmnVrJCNVodusfT
TkkDVFAaoDpyvTSqDhoDDuWlmsgKksV8GmhRbyqus4CCpszx8Q5gxwaXF87frXvb
WpKVDKCXWBxf87bY29Niun1HGyRJCrGPQsbE5K0aZGx6X7RuxZIJTRjdqFLJjK9E
ju5QWs51eT7w99OPCiamyEmnOtfMeDSztvtaksGJZ3j/9021HlCdjwd5gj5nhgOY
w11xOTszpIEMK28kw959PH3KDk0Ut39rudVMIDbR2EfBc4lz6Wkzoz6ygTswUluC
ccOMFXBmIv1Go5m+/yzJFo0UnGdZKKWYROSl7CPsMZcR5QPYEpKJ2HbyB2UIxxMK
0pcwl6DnkPQlqM0j6ipMXe7Am5cjdxhIni8x6BVpNaUqXIHk1MB3BwR6B8sqbVdY
FLKR558GbrusaYnRY4+YqEs7tjnPuzRLzqMZ8H7ImCqSqPLrWXl3NYQPculeJPip
3F4DQC/XUwuFdoHgo55k4l0yuo16/EPhs5XTfUi0oa3BdulLxcilCp+k6c3dhjxg
i5q4NGRowGBcNpKNBQonJJ4E1tnlCRMfzGYWuqUkhQ9MGXk1NugPPXWZm4ijpMlM
57rSjufMYNLg/qCPmpmQ244x884ZmU/YKFfQ7b22dh2NSpWobadIjo5Qy9QOHSma
xS4WtyQ1paPTay9QsPP22fM31VktvB6fMZiMor1JnuPOObmOjBjyjA8DbVWMAjgS
czZQo61c4BPsvfo7PigZgyMcFxTKJZRSSihSEPoEm1ChFyZjgKbP6iEFhZDhMytz
ErkzJOmIKkUMQkt++lxcv5V6euLh+/8HjEuShNVFaHKs21z4NHnWd4U8ubEbdSBw
aN0G4npzmP3tYogYgbqVCxFHSNuMVwLv5H+E2owx0OkdLE7g5vMx4fwRBpR0Eghk
f0s1qZiALgJxKnhSw1blaoDbruvxgGyVJJG9lQdSfWpnY25SwL8VVaQHa/o+7WgE
A1ibGAJ2ctalFuUqQVUSg4nHBKlACkujyhU0F+Hut3l579yFrlejnrMQYszvzhIg
463VB8tP83qnvXLx1XhU8mxEUA05QFHhNTUo4/m8RVBnW4W0q1de/xXkriWuE4jJ
jghSOlwQY8odXz2atSQyb+PlIGnHC2cvZfRIvPiwGU1hsVTVkn+rMh1DHRQvZkgX
PnMXPzhk5iG/M1zQNhPqV+MovQjS8+sH5zvAi8SwwT+mzWNAxIruhir0ZqUO/so5
+/o5fGn68YOTy6EGZGD1X18BaAFAASFNE88pd7V3A0vl2Acb+U7k84snTni0f0Qr
h6iVn6uqIsdKjySHRQ6gR5iRkVhUUwig8WhA10xLDu0MyliI8fBNpJEjqXSUsA6s
uav7I0KGGqgpd/GMogXCp49DVil9Tvid7kWy3S0x5k5ZUjQddMHluzSUB55BXTa6
o10nfQu/xpN43WoVi2gP44bzfj+sj3XVqqgmKvNyr3uzZxfrvI2TWijTsKWA+tEA
QEYM7cdY0M+tR55pWcJwwvFpa9niKZxLsaj1IMA1LFhyj4Ys4k2uzzmBB1efTnzR
wVZnjHY3FnrxtgSTvkw+7fPdM6oQJrDcq6UEROLpu0sYjqDgAM6D9LSxkQgzyVQ7
37WxDYExGdSsD7WvW+iFxV9OkvZaDHKVG+gf775ZrAsqkrNz1xYvaT6n5TC7irtK
LmnCIg+fEUYQBA8Yb+BEWkz/d9ov2mUVH7phgQ6cG+js25fHIyDzx+VgMlrJbYoH
OAZ62Wis225MSRuNBF1/IVIaa8USPo/geMrQ4THiFrDdW44knorSB3m9Z9PQBWj3
5pYUIgDpmPZdHeBdG0BM0y18s9NZCArDvxMfVHVdZdqncXpK1HWISo3MgVHYQDxE
kfYlfDaYAILdmk0M2pvrlypA8K2VvYKf9mWAV7xlHrpJ1tTSYDlFYewk5YELmXuL
0z+7NL0Ue064lZ7iofWuW0QaYu/6fPrs0oklho9qZZV/TNOYkXZ/tE+8F0b824Jc
rTKLz4WwLMuTvrIUmDg6zZI3VUDDSWNMYGvXY554wuk6L/+qiIp/k33K4dkgS63H
MBD2PBhCTeDjqNbfawZAkq0VLxP6C7RQPQOmeaY1NS/5j69MzN14S3hjByFDEBzi
rb3PuS34yWIB0dRm+YZCKdXUuShCbcK9P1zILrQHj6Pz95timyrW42aZ5z/KOu32
/3cMiQdrk7tEfmHq5ghJxm/bRq1CJwssPbVtOHDg3TMePVhCWlaMgAhhjuEdswMz
rTnopiln1o/Z+mv+Q0yIvcJfV1KHGMuhHEgRdKbdqRHXylASnRlBcZWusQml/dAi
cH/vLZoL87y8O58v+4kDycNHf6nsZP5ewOS8Vm2U/BgXToIaRj+M2Mpi0HgEcBvn
S5PUjvgkDqBqsBcN1gOQWArQS1m/RMRPoxmZQNMYIMIjetcwA8FjDKrZmw7Rup8p
8xQE5ILfbhshi8r/PGpeRCeLrJMzcGyMGFFkdyR3rulyzaCpNv9m3F5ivOlFdm5O
lEc0aod6MWAViK6a4MZHhmKvWbVOUtcmY86ekIAf7jcS212+kReH1HMlF//kULNR
YErivPRJpGjDpBRp8eMyxRiCHUpdKqMUjDRlGraK4Zuk0GYVkyW6MFdMf1GHOJAI
nZhJgNlE9vBB75BYFERpuaVGacMHBxkZhm5iO+SMU/TJUZUL95xFIP38+lfy31BX
rH8qSfO1lpZcyL9gbJMl/SiBGOl4cV81BsKykCITBHTSJEWCm6xPMvWjft0HUEi7
jeHK9Tzu8nKNTPqRx/Lqq46NLz2xDSgHvPJrIIh9qY+wPL1s952Qj8hAKk/eJ6SX
1DY7bJlKFUgV1x2GpPmbDJVqvZHHFmHvXaYvtimLETWd7bNCsfLN2gcWYFrnrent
DPRYAfNyMiHkQ2bLJh+uf40RH9nAxBCg7qJZKUnz0TKKhCZeF918EWAjTDj0rv3l
0Zxh6e+NSXCallcEQL2V1IX+BeouTw60vBsDOPWWEWpH+NqaFwwfZPPZh0BqN7o1
wtTdehOdh1AVzlG0YefKLA0SHprR/3Dim7iNerABPFZysN3LKAIStMlnbGGJ6jze
axBBg3yUUG/HTh/P7MIzolWYtiM/3EdWkA+j92qi58B3kZP3f91MNje98GNcooPI
HHgfil2FZJVs1OvIYeGY5z8AMFc28Ff3wg6vyvOrM06usJVUo90t8UGG1Ln/R3f2
FPbVGVA/7OkNOKq/6QpeHh/aKpJGAFwige8Fc/zDYRX9n25kzdFTYYyvLAKNRfWc
Xa6l4c6F8BDmnquSshpEiptk9g2ditgpU6G6YdGczB5rT2bxW0Mp47ELeJDxVEKX
umBL2Coq8uXMSl+meeyEHIs93MGd4odTvZ7dLT0fYgou6XhJkNp9zRFpqtp20NLN
x0zSeliomqihqcm80rBjkOHzk5Wwlbc5zW0pfYgV7WH51wGVPTxfZoniAuNSY6Tq
QD7WZKKBW1sxgNwVaqOggh0HK9Ivq9qsUonA183hjP4IJAeR0syi/nXeXoRHFpBn
V+6HTofMTiQdDwfkD6Hzz2ABgItqjojxRlBNrqj4WKLcyvwpnFgBknnymSyHMfJh
4G2/4nvtLLX/h69P9DQ91RPc5sSbqIGkDoXaeQSSXLEGeci9rUKrJnjkLPgSS9IN
IHtAqESKt4qFpXse2GxmOTEJd3T3ci2EaQDchVNX6R3rtKTYnYo/U5zONoua9yY7
5HrFfl6EyUELxSce+enjIQfu9raMwxQk6QwjAx+e0HAIRZyukAui5RO8LaySLQCF
AKKPrEMVwYhcJDEqI5rreWGMDeqzSmozYIZawOha9f2Y9m/TSZK8Tuz2/930Xl/Q
FZ6SK0FMN0MkYhXFXJfqwGQLA0ekXcWetWIX2oIyb6FiCg03/3ByxqIgUuj8kNB7
z6PyHHlJj/kmE2TwOpg7dSrYy80CC6nuQ3qjbOG1czBa/b46I8UCe2DdBJ8K540B
SEzvVv20Ki4DIZeWhks2y2/uU3wAvZRzZYJnZiG25h7ICk4DCY0M4S6Czrc/R1ll
ph2GlbC4ObiDItilpqSS3Ooytv3MbAruvd1UECOY/RW2JCNM731YbPQxwV/BklIg
BmzqbPL1O5IgqRpTxbZyRGbM1m6BSHeQf5dkEsWgAbPhlMvFRf4aggcgROOqbg6V
Q4yOZGdlMNWeI5w0XB2NbasegAhe9UFZNp8hlmW6CFVjR/RQPVRZy19b9hk16Sj0
5/1su8YAmSonzGg4Gpg06ThQK2y0BHmuibC9k2INJUkaPET3qRuLqtD45QmCFWQd
gBZPR+RiplmijHuMZOb2e1FHvYDOVxI9HJs+3OHysO6GOtx3UqT+LUy0a1hj+YNL
Y1xums0FU6LjhCC8bRYqy1GZSzgELylDbV4G2i3wFfE3D/8MJ69zpFQcYU+9vBYS
Rmwi3lCvwCQQc+ILJNsmRKCyZq2n/ohm7UrLNSx2mV/aGjSleGtznkkNrhEwSvew
ZQLdSAvLwEAdDtXnePpV/DfWluIP74BnWFzbM6u/vkUwW4JVams5dJntEKxH71+a
elEhGCz68B7o5TgRyxoeJdwFGzAhK9dmDbygXnUk7EdVqa6FHCXd3RQF/sKWmR1J
Jhthr32IX3USgv6aw3t1IeSIQtz866s3POxMj9O0wJCakwGNCY0Wslg8Aomgb5hy
stX+fzDSFQPyhjSSUndA5TQXfiZVHfF+yRzP0tskA6ucIS3rt+Qukj+tGyCVvqaB
k88sAbsbf4Ex2BujPRFZArDKHzIBNlaRUKs1JZP7Vn+A2u8iXKwwux+kMWOs3HvU
TaL7fJCouVIA8+Rg38ZSpld2mEhsGfdjELRmexwfHm2A6lV/alze3PlwSSm/BJvp
inpVKB9My3/t7udy9fUdMpSpqkqjkMGaNEWoHZP/q0cQzqYf1Lhy0UjNH54UolBO
WlUvS6FQaS/zUrPlLVxHB32K/BhXfKuxSM0Cy70In27jRF2NiYUd1QsHxs6WW6dm
24kZoUwU2TtrXdC+d5z9/nUyQJIqhfjx6h31x1qE9cq/eZiSaDPkxRH/VJ1pVNww
wOHBw9T9HsO983+tfAcjuTdWbftZP9sGrAjeBX5vTx/ztZWlK4MdM7Za1jCPrzv0
1Htf/znTGlyda90O3kNAHswOZelgEQS3Aw5UqbkBQS/U+SlrIv11hC9XKm4gMcLh
8lH9BjFZTdPtt3XjnMXzDTtVeI2uMU64odDsogq6wADcBECTgoICMJxzICrec6o0
m+HH+1mwqYafmbcXQUzZdzLgY+Ugn01bIVN8Ic7vrV9hhNvwzszCwzSHGnThIeXg
wd+07w/qAPk8i6u8lkbGnSAAZdCM/uBc1o/KRurUSiMxudB0qkAqhA3L7lti+WTx
kGUIEiBVijIwPis38Dh/diQlyIrN/J41vUC7z2BOdh9Wn1E4s0SJdNliLnMJeM05
WqmJL+Wl4ZeQcTCdAzKnn2G0ZKwDCBiLfGw3ehShxTlh+yrpWagugcxApfd5QiPu
N7UcUAe1wpACeUdMvKNHPYeaGFR8r6JOUL9vI5vV7tszlR2bbUtlDgrbCFAL2+Av
SQQCKNuYHAeAojb4Dj2PMwmjpGYzQCPRFZ3sYGHGKpKSAAnLLrxjo6OWXj69oQ/1
y2PBv/CBMnjtdpfvVfpoBb+2ff7kCOXue4KoA28GYjKwwwvj7TI5muRN9aO9esAq
xrodYKSJ3GPNJB7u8ory1Htb+3aRj9f1ZX/B0TtINkryTOAdKidWqWMv1UhmA7fN
OU6UZEqlh+473gzym2HpfnmEdFQTiJdKiVaPx/UWaA/tql2OapQoMVLWQEsCV1AO
nrHJtlp0sPsaioQ0s1jPkSMb51SYQ3EojUgy7HAOJYKrylfZIOYFhohrdBu3RMmB
mr50gCDlsyFfqlA5iG04zf/rvYP4P4BI3oydFyZt2vbBoSMH3/jTj+IGOY+bAjc4
md5bk8IjiJAG9Ha+3i5lbDQoIKff16PUUfAuB9ouG1PLLljjy8D14M1oj5QqQWwy
gxUWz+VqsaQNRS+OjmYHiac5IqVLoChESrq8FPh2wWxoyLA2U06lNTIzL1SiMU90
RH5r0eeVAl6GtNfAdXqBuT5nWXAi53B/vRFya4OxG5C/J28UJQilUNwxWAvsa5vT
XpANguFxRxpPyTHTUcYACmYkDlflGlr+h6YFwLJG2rxNepaM9UXgXtnf+73vluzF
lLwCtoqdb47DmHia32P+IbV5J/q1KhwYibU3L6z7QDekC9m2IkzrZhj0sfFQy8fu
9acnMt+L4AH39+gLwLJL+c34r26NFNmTCuqtsk1QWbSgcaQyXOE+1qp2G9x1TW9e
6gJyLYg+diEl8FIZqpWUi4m8Y1Ur5A3x0kfUJSdUeNWeoeJbz21bq3zyf69E+Iov
rzbQCwRPWdK37Xv6oWV7PTa75hnlvZxIlp4n6idrNTnk24TdMEdC50JMLrvJWhv+
tEeMq6BRY6YMbPBfigZHwx/gN45rd+wOyhFFs34vqAWIDWfE6D4FiNlDBfxpC+zT
SwNPf6HLdpcG/+PNwswgTPjr+idoOp37V9geu/QILspQ8BTvexN+MSv2EJlmbxn/
WE31q6FrNqB5rOw5Rwfy4D9wMJClhykCySzn6Ck2Ps9cwweyaka7V8u5sz7KoabO
xizgEmQWZ2czqiGfklEaxn4RTW1gvT111vh9fNDfR3ahC/UFl6THS/fB2jUJ6E4+
bBmpZyxyQ1JAhRhYZKGKw5veXCTzsUCOO3faTxd9T0fgUc0RGt0nZ4p+xUziodFT
Qz6iTuTnrUxGNWDGrlbUSjdztYFgXpExfuLzhDjpQ7hTKl18oEKxtZqZZe4rglsO
IpnhuCZvW/XzjjIFIZtcCQ4h66spTEQZ81qB80qct3HXVDQ9mGXdgjFSu/ccy/T0
LzBKynjZtSfxZ+FXXtER3psnOS9Q8ycOJZ6ZVgYLh/hYkq0Ilt6GSDETtDnJd0oU
QuC3IDC2JOH49MYfyXLJ9tk9G+IESkBra20b6AZK0JB0rT4RtHRZ3XeehvwzMq77
0bsQZMvU/HiCeSbNastGP4bOf/fGwJl9we9xfxBqaFyXM6Cq0eOn+uuD7SaYJWEM
9Vy+mh6xIiYFBPxUIrvQO4yiMGQm5eqRkTD28Dsf03w=
//pragma protect end_data_block
//pragma protect digest_block
YBtUz3zpuigdpfr5kxcE2lpj6I4=
//pragma protect end_digest_block
//pragma protect end_protected
