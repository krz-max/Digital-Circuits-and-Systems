//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ANc58LGfQmQs3dWBuUqqgnYBNAsL1gJlR0YpVc0z9xv8KLYLvTETbu2ufZJX8Vh6
rNdivhgpBzTvD+LvzUh+LQLIvFt/pubEKscS+xYOjUuCHNfkWdI0xX3qc6+gQ4ub
S/x4WBpX4lUg8xEe5Smzntk+kNR3T6GyK3kSLY0ENhZgDKfQkyk4Yw==
//pragma protect end_key_block
//pragma protect digest_block
g6WAfmXaRjOcvzIth6zt6qZx38E=
//pragma protect end_digest_block
//pragma protect data_block
OkFIjZrXFEte+gBfupjHKiK78caC/9YYplUz2JkBGZYdqugCHl6Yhjl/U6+fgNYJ
1FtZUAGD2P0lrElNG9KcUVUlJPNrjZW9Of5OZY114/L4z39zuntJg9KQZBb58h+u
ooyQ4WJ/saeTKpP/5rP4t3P02T0wvj0FR3qkjbnjuA53YOL3EGRW1hxbrac8qAF3
WEZYK4VBelCyeoFIy9Mxdjxe0dxJL6T7pR1LZkDQ5pIJ7RHPv43F5dZYRAEkr7Wf
uqjVNs98+i0M81jvCNhTUiRjCo8L5GnqNGsDdYwKXHpKfM71lNjwdXAnvspENh42
FCY8iT2BKkjO7Zma9J4yLcczP2gA9EOpJqhMFWv6bguk9kWvAGK/2XludoNGr0UM
Nsib3/ZAw2lFf+5TwhsbQsvcTHmt2kqm9RL9752SGBaUs0jMSP/Kmn1GaE/Jsi00
mt3fhEYKv4hbgq1rjvJibcxpWFbLlvYYR3GcOhkL/+lSjF3pjqjwerzkK8eT8kYm
6Dp7/DYG3GpvKdzDCgPsy3BgUt6RJRdVMrFHvQcWzSP15D00Rrjcn7XYWqgiqDTn
EZ6xCaSaiM4c5NAJoD2V7jQ7qKIqt136HjVdPAd1iNj2JxT2HK1TXIW4C0Ia4XbW
FW5cRGgO61kTx8HzDoPdarE7nwvoKh5u+8MfJK7KaJ/P/OvxGnHdJSF+R/8fi9Fa
h8AEf3Sh1dOLr9YcDwXTfKXX6YGCCgvNPJC3Dx3+gp7d2Iy4ADhMsTRUnyQ5/pkX
+iwLFJGTkM6thGP4Wu5tnO+ZRYzKUnBuR8hO5UtoOJnI8/lBzx+Knh9TGTHO3h+R
mWCS4k3Kd5sS5mYHQUSbdsJicECyn/6fuOWBlJHVcaE9F4dnFoMN9347rKL33LAi
JtUSB6LE88rWGDMl32i0eP6ko3DJQuJNy9WGb998jDD0YwXc2IQj7TRn5Lh6+zwW
Qm6KnLJyqJ+DBCHWBXI0jr1z/8B0bdQjuiKERkqnCGWBaiBif1KUOAhuLoE26EfC
Gzer8Dnd3BpPiVs+XEVAxRqUPwtYauPDApk2dxYOzoci0HrETpbt4ZipptNAbatn
TRV8cxfyboDedBok2IZqgxBrOltncrf5+0nbGSUOGyO0bbk6hAG4IfK6w0pHkEfh
0TwQOuMe6UD1Hoedg/UwosQlj04VkF9LidHqmXShDoZXeuQRav7wuty+8/W5uQKQ
XYRY6TRDePT7BITfrLkSSibg190oT8T3xX6LlLSQlOgFEFduqBYUjaL0vEuY4SSI
qgZuSbisB/+6Kykufqk1baUXW2WaJ/I1JCwP/vGY9ZcZ/GMf6RGDAf0yd++3woyM
BZh3bnpqQfWpb7FUwzWLmhhBck64cWV+BjxH3GOeq21JjJAjzu+uo8sTcs3pn+3e
ZZhoDP7WTKUDBE3if2fRCbcFMLAh4WZTrHMOiOQQa56JEZhaiX+uE38G2DKZyJMr
0FampkKUOm8NhZoPWuHLC+YuCMbtUYv1r/gr6glsLArHkMVxV0Jqj1GW+Em3Si2u
JgHsfzYZd+N4ddmNebqwUxa8MSyaWEjCaEPY/9EDpPPIGaTuX6P3+xgCX89BgA0K
3LORKX8ceLCLmpZ8eyyA7NJXu7vBCqrpM4gPjkfqVXLFw1LAqtiQovgaIChwYTqL
IKSAEwKIu4nrQIGB3BYGLdhhI6F1LhZzdYE12Y7wRoC5unPhbt3IfhbiSCHKq3jp
QCw56SWPBDjuU3q2FvHR3o06kIRfvGcPrkc41gV3f2/2uJl+DbxO1OOEMCJqE0II
1eHQrLxP626gmLIWdDWZ9OymREU+XktMDh9nhRzd1x67ns+HGrKpDQ7DM924Eafu
w1CoUQyBf0bcUmoa42KXHO/fDay8r9hZ2qboHOfLhK52qGaLTHjC2hSUz8VhsUbk
IPWf0dY/kkAEELRwtBc+JvZmUQOiDSerk7Q5KQx+MHyktFQI5F5/BabkJ28jCzV+
oHB+7f7xS9CsQS+k20+dzYe8g624xfglvlJxbGXOZeUdQItZ86M1O6HSxGwkv47H
ZrceIMaZ/np7J8TEcGl0tXwo7hx24/AVAbctohel/ngsmq+M2S2LPWZG03MYrmYZ
jL+CRDmafClozepJmGxd9gtPGdHqF4VB1BO28ZO/P5SAeSvK6kJJZP3YnWKFb3rO
o3yGMIhNCmTuZ22pgVdxTjdvv0KzVpcKYp7bVT/P9IMggtd3s3MI4i7VsSrdxoli
oTwEwp0mijYSQzF1gSGNvR6c2oYpc2He9db93ZG1s4pdPXyDKvroe7Ai0oY2UySO
ZXNj4JfexDlyIcHVu55HObAKBg6TWv2oSFHtZ6nVWZGoAP9EkDUagTutB4OVNPmO
2zD/3uTLnpuTJJsVbfIZdq+oP+VcTDhXyBd5w3g56APem1ZG2xy0hKJ6gIVPgOyl
W0rvpXSAAOMITQFPTsukYdXPVXPJIEY/xC0o+cd7zCMeStfExBDV8w/9DhVF0ICj
jsG2cfBcLu+zPsvi+iCdksLgqAyWZ77vCFQK9CsORGy6d/XI+kPcMehqetCs6zlu
iVFFJgNAE2hpxpfkwJSdBcG8IhLLmluJ2fLVfs3Z0sKOg5ds8O9CjAWiLi3BZIo0
IuueJ5+UdoLThoHQ4ZWbozTU6snqTmo0ZfPdnoSkXC8r8FPxNLWKEhMZ4ypfSJjY
+BTn5NWgps8qFJoZ9SPVj9VoCZG+v/x8oUl2tr8b3Xb0yPjyRLB7VeSa1lu3uwrV
mzk4ey8p5bdpXzSf7WXiPyVReArs8LtkYtx3+xAKqQVYWX33TgOwmun0tATFrBuf
q+YV7yr5qLf5PhP95MBxHzFg0oIIGmiLDUwQKTe0lmoQGPbsLxK9lDTpZIxeRJf4
eLLY8vVdHOcmtw7dBs6nYBn7J7bgyDxaXbJj3ObFSfQ8tWvWjRpwu7E8+aGSyB2y
rZRoANU3EpHnv/l/k7VgNikC6+O4BkTjtWurBJG8LOHT04e+2ctnaUfjC0yuvK6n
rvHS7mVXyOvpFJLTyGmLKbecvuyWWAzVezFT29XA0wV3d7xy2P4LGXxsjLOEg9IW
LGvuEnVk7vgA8K2Ojg6dPQ2mOQAaGKooo3uxpeb7UyCRVJRFPOBqGIE6Xu3p3v+K
juHUav+UWBDreWA1b6i6UKsqoPi0OhT7lm+yoLFDscSo7JyF3EpYbxkL1/5vTEts
uR6SsC+PiwWkXDARn3NNogH/Glj6NuaAQy9CHqvbUeIQcCLhJE8UIfoCXN7c90NB
HHtmI5gtzEySM5KRi4nTGOitjw8YTvbD/4LD+BXKUZL08rRtL2ckVDVYH4NtzU6B
eKO1ZhC/zVNXRbQqBSFyh584puPl7o5zNplnZTiXbflMjAAg1hJ0A7RY82SiLbeL
Qom54CvWuWJcI2zBOSs9isy5DI6eGKtVfQnHHRCY8p/CUMIgwtfHma1YN2Ab9IZe
ZQAcnyTSCJyvMj7rV+Kudxw+VdcN9dZpXMbzvnj7GQOxkNDg44nTXmHCpBVMSpxJ
fQvTl2o2GdUSFSrFrVvA3X5QHt3dwU4tDe1oTIvBqS2spCIf8nvelHx/nPd9BBy+
hKAvGE+MGCJOa0wa2uUx8GLkpBd/lhCVicOslTjTnx+O0wbZXFDaImbwi69gxeJf
9lBXzjKsPGenL3HyvII0RpSvXzhQk7YuSXylUOoGQhDjVeaPPAINZVVHLi2xZpdr
+pCcL7q45GtKNWk+JJ/CQREE4/mneDGRsnoiJzJW1jaFvrfaQXxINJtz3nRx9528
ITTF9QIbmbC1tEPkg3ZVZb8CDEZXrpno1JTkwBbfAj04Fod2MhBahRPNcU+K8evy
p/GMB7lA2s235NShYSdbKic/4E8E2RJ1l+PEv4ksHB2hchrUL1t94fKqd9m97ytX
aTttmsZBwKoOCNxZWEibL0moujK4AqaSiTpaqW6R8PXoCvnsJeVzci1MzF24pUEk
pKjlDl4Yn8Lrio5rEVI/x2sdv9Ak5MK+PTI1uioTw/7efidgTreTaBVSqEQz36cu
ADMh9hC922v0zGSz1ZYLr/SuM6y251vcJXKeIo2pGXskhAiHNTJo4NRe/TD38s2z
Ln+4qjbpWcT5qn1i+hr7daXaMx2zW7nm3rETVWdv1KZTmSfQrWfea+gW4qZXOOkB
EqP2CsfS7wIAh+tKanaxHDGRjSxzAkDLbRAAS3DqrhlRlhOAXX4TYfGs7o3EJ95U
8h6YMBMjeSBet6WHEn/f1Uk5BT82zMPp1/zCVKLAsxa/evolDdvlyUK+fl+y/u25
EzPyM9nAnS0rjAWBd0T6n3+gsCjYKxxs3TJKwl6KgfQPvyIT1H/1LME2M93l4X+4
yzwfiG2fLw5jiYjYk0F/7HVZKVA7/J7hkOIWmY/5OD3xzGghZic1Oklv8IlgnbX3
gyC776FLUqoiqwc3ZD+wb/YGrb2MMWrqrM6U+3EMh/M0R6GiNesB11/5fXpCBrFG
LrffmaFIo1OBE/uIDsPIJNrzGpwdMLunBr9oVYvcZRH3g1tCkt0RjJdzT643EHU6
jhp6h1GiLuYAZGyWx/DO/ZIOwdcOZecyznkz10Zl25A9UA+YcEX1FVMQRHDzhKUe
ImLbmP3qYGnAGxLb9tDz4jfFJ8CmY/FxU65TOf2HTT97kBNwg+q4UV1+dWM/sIuU
0xuSFOpwZG3yaWQZ6/Q7nGN+8DdjF+XV/k/mhDiT48SEXOr8tv6+PSstDsvKVGoT
6vMdiBz1pqdHtH5WOHWVNWaqsmvO9cD6/5rlcotWEV6WtJjekPDeuKvbPUpzhrXh
2uK04+d8a99NALboOKyTXt2Zg3IPpRzLDdhAXvWdYM7lKNSZyUNAd9qbc7CJksRR
tYyo6lwDEAC/0Gv5rBQQGgkXNNevz4EU12fgK8yBeLJM/w7Z9FtmMXfU6dSkK3me
qsgv4CyQOmf5ssCsJzxrtz2PGM5I6higpQrNAryxgBMOelCwv17iO9A2lONm2cAh
v2Jyg3jXJ4E5sXaY+xyP6uuwxKR27j8WeBuylgL5p5XAgeEtSDvwc8hY2p5uC+zJ
PHaPKoPJBW5lxMQF/9XvlHgpHsUrgHfUdjG4qhDH4GMEQSDmRuhlSkFQNEgLbPv+
5c5+Oqib9ojRxUCnSnXliGtwbhRyPsMmjrHyEStovjqoZc/PLodYCh0OlPzGcN/7
29GvF5JmyioF4VvLlV0vvSh0FKwbBt1J3RsowhsR1B3iD3ahNa43aR5f3F+W6fpM
GZ7ZlraOm8idysmUz1KMoHNfxd+eD3+xk6gryJuQ7aW2qtTuB/cbnJhhzJweQgrO
buEHby0gG/kbDkBN+g1mTbRYO3l+gjXXdV5IGf+CC2Wuf1c/jL/KBOQMItPdlJOu
ofD+eezU3JnNjor7LGggd9YM3GJgQMi6ajGn5OsYuwNy/RQY6zToaOOLrAiWSAym
fKqrZTlXtt0/yVjhdP4vzGx7mCFMtQ2TmNnRD9e60OoRk+OwwCj613mGek+FEaJV
48+gn+tBMTuL+gukI2g0ER06ikaWcSCwK4J5yVYc++GtuGYT1VgAItnGN98LkCCf
m9IFVaD5XgcDFMzvVuVEB0u1kuyO2qxZi61U7R8xcBk0eWmb4rfAu5HAhlkMyx44
SaoAq4J/d+oUKsu6J+GJnQx2QaTM+0F271OHBmzAFtktG2JKHaVmVZ8Vp/GlyRLV
ChETi1CzEpo97eyJq17YUJxKLVJxODrXqcFb77JOM7uIg6l+N8uB9rw/ibF/j8sM
OG35uwfdlC51BmsvzuO/CglNDTwhuWvjr4CeRP35zfgHupZdoMpOtmOWfqNZ9gq9
by1lSlHXC5zoVXQ52EktfGukUmJ22xGZPDNvqTlyW4mpeYVe05R+W7mrMzrC19WZ
Bsxxc80RJwgRuGSCBI+4x8JcsaNFZj1KKYxmyNU5MbeDqeuulFT+o9vafrza3quW
yNMUH9v8y40P0xg5miQSIFVKvs3/V7SiZ9rauFD8sQ/t1fxx9bsoo/gPeABcBLga
HfKKH0fDjFb0PvEz3JiA/q7qlYd5JAQZ5aIznbGH2QIaOSM6g1v/xzmmytVVq3rw
oScEvcrq/kkV5tc5mUk+1zfZBhH4CK6sHc39WjUkbKUBpbwCvGYGdC+hHmOe/vZL
RtdxrKJ3ElQbHM/HLWHlzWInTV8MBH4ssZevfuXffrdbrlkoErMh7pe9XZiqkeoh
/7f3zybpNUNsC2KGsbrTd3TBpDLHxkU4I5Q9gQ5+ALaVsI7YnsUg39XB1AdC6EAz
dzvS9OD73A+lvk6IPL3XwxzKGUS+PS84oxI94Z5oSSJS2y4P/OjwR7uQvWl9cHjL
a6sGjE/i93bj9yQee1JfJvSQ8htLIF1oVn57e1bKTy2j+h0s950y7OuB1RkHsxZH
4rsDGnjnaB1VO9zjCJTitPJ8j53iw+xMwtjj+zDrM+Y2Nm6ECssaARtdMF7FxjBC
OZSx409aQpUGcb9KGX14kVZHZxBVirbi2C2k+B8WWbxTzB0fpUfe4ZRFHKV/TQDX
1V4qV4j1oBiJ3zcTPk3NOXbxfANCmhONvbpPDrEbct5SKOohaGmnZ9+NderHb6nQ
215oEBges2S4W6dzKBOBJ0VqgCyahmMKtknfndkfB0OByFUgpmzsnNVc8Y112Cyw
20RWFtOPhDcSswz/LNfPd3eSRS8rgk94gzih/OwvZrR3OJlQw/s7JfgxUvimet7R
p0ebycMZORP90NvtQlEpJCcbyN2Dbtc4NT8/KRsyp8av4J0HRcmNViNtF17HCGtf
Sf07HX7qO4/U8oTIiF3Qb5DI0DIlVtjdyCs8DJ3nNJBmSbo85Cx3DkMTz4pl3GHd
Z9k+io4hRkpWAGfiP33AQOlYDWOJPOrRhuc9w51D5o+nKFo3KKszjd9pK81HodPz
8qisgRlEAmPsMnnhFaZEHD05PcShUQw4AKFScE5FvO73DdWyQ5ht65wVAgExq+pU
rjd89iIkz6XmpGklHCJVJOJb8L19BAWX10FRtYHzITza3GGNWXRMeufLyxBm1b4p
P+4ZEhlEfpJhvRDnGdCppM/zbFtgFef4ECBbyfxXiuKO/qj2mZQ7F0i5ooNigXr7
rwF2kay8WG9CDKfiiHGWlculzbcyIg2zjaEQs1DBImvZLPb9wLm0w78TzZ3DgJQz
f0LtfMbwmQcAUNLkURH/RadN/oa6SNpTqmHJzbILtgmE5DZZ8gnJhrKwa7Fzew9d
5Y2BZvbPkxfMkkJrIuVVwhkUUqF99kitDHgZ1awSqhI=
//pragma protect end_data_block
//pragma protect digest_block
JaO+OliCL0ec9KDtczScN6RUqaw=
//pragma protect end_digest_block
//pragma protect end_protected
