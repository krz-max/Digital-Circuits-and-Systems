//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
zMdDObFJhgwv9vlPRm2KPidm45iX+HIH+IFB4WzwFqty8VQGf6X02/NDAzfiq7v9
AnZFN2VoJVCq8/IM7oJ1VzZzajV706vgwNaAY+dKpsbsSmOKa17SahIxbeO8vHnx
80iTEq5g36FTJk4l2fLeJpAB/y3EDnBUDDqnJdLzcj4+ufKL44idJQ==
//pragma protect end_key_block
//pragma protect digest_block
G8rlVoaWbs2nGRksMTZIOkmIjik=
//pragma protect end_digest_block
//pragma protect data_block
m/QD3LYKTz4zxdyu/JKoK/ZnbN5z4iwGFgjrc6EkTAyDJbKy5BDbjeRegHlijnvW
o1viZSscaZmQFD17i3Q9Dx2M/YlY2qFjCg++6S4Qf3S5+sWrOffZz20zn9wSj32w
54Yk/5bnyLbwyVZ1+VUCgQxXT1R3g/Wf4SlBXerjUal33bDI1JJnL8p82QZ3XsPd
URdqKe0utmisl8T7/+JldQfFjHLOO4JLRQiuUGBhfrnIt95l3QRXFK93rBiIVL0b
vqgczrw26Vjmvw+zil++VDY2WffgK40MNrd1zdy535/J2VAC0pxSeFdgY5ZSft1Y
/gIPtAnLswqU46UWDYad0Cp+V1vMEjA7tqBdSD8M6RlA6p7io1VRInWTVkA9s24K
RyZJdtFfRBs6Vg0adkXnozmBrXkOrQbQs95MuBFKxQBDXWjIBuAAvwL/eSMei8n5
dd0lClW0mZeTxx543gMEP/8oNieH/z4nAtLTNEkdmTpEwT8HEMvCfaSq3VCwfQ07
GLgt6ag9aWc3yJu71mE4SPsF1KGgNcu08wWm9V+xK02jaZ3UNohEQ4KbJvsXUJKx
xVrl92siq/qpJZ3ZRYZfGwdK5MiN5EC4+FFEa4rfx8ZdoMHRVbIo4vPH4Ay/T1yD
eRaKPhKloVZExTUHij/++ZQV5V9JjSrYuE1eYcDYsshJhY1RrHFZGmCaUIloIuLQ
ZqQrMpemrts4yPMm7PzYmG0R0l3KoKrSjmUNV7qxrJ/M9cCbYsJLSiPvEjrmrahp
+9Gpef4lSX/I3jD4ao9i/urk//0dz6TEKZvBip0Ir+K9EgbJoeUseWfzI5JyLG6/
px0V0KgtYfsgQXRy7N3NkiArDeBNhDwLZq6fBWIqGBh0drSVZSFUIil5GtMkaC+S
/7+9d4tlF7b8Jy0j/zNUqta/CWt20r71IQ7S5x3hmj6zvXt5LNYK4v3ALeeSr88p
KtkEg1/9wfNSVn8CEtjTMVBFSkBGkbBc+vOA9oh16DcgvXifgETyV3Rc2qo+4HmK
VLPYXqoeR3fAgWjdFG0mOE99uCMbOVA7nQ8vVolIQ1q3FLhfKGde0V6BGzQiN5TT
PopDlkGAibXwHETUBCMXbn29kieTEdxmdVi248YaC+h9tYizZq1HM6KEVkzos/8a
mbuy0G+YqsVHc/uBUvoKiE+86O0viRqFMZ985mqcd0ivuJsFOh8yhHrfmGNwR2k1
SO8N39Cng1vOD9DjNVFs6HCcrbW3B0DzpiKJkSJ/gd4RwdLmttTFrsPAi1162sbP
gp31QbKPuD/6BQMWnWWJ/2onpoH4q7/+acu4QUG/4UxZUkTXa8a33qvs1shiZRUb
6E1qAegyfxlYAa4qODaSTnY0+2mQQ3RmsOO2JrBY2qiQOZwujtxrFmOLM7bG3+JL
O+sWsGq4qINIW17UzL9/9NNy2pCq0Wez2tiVF8D7HeVgObZfTg1E4ijmoCp0FeVR
f5JP+jzPlZO9E3V/+p/pFk2BVVBTYcuw3AjvziLs7JVJO/7CIyDYSi/yODFF8Vcq
4QraFhQs7+BsNsUatbJMTjEfqa85H+a10jEmroFwbrlaK4xwDI2RMgcNtqKK2dFF
/M/cf9ANMCaNT4pudoh7GuNru/DwNckt+JAsWIqZl+g1SCYp3e0R1U+8YSDCvrGj
QMOpX8MwI2o3wNryh+1z5tGoTzq2u5iiRvGGtzk7Vf38P4xsDFX2saim2aRZ2nvF
gCfUDCSP89ZeoOG0sNOnWxlY/1E0f4htyKUxk1SBUSGY9Dk3TLSiNUoiuOEzDZFY
9l8ZHQYLS3yigQBjdMDHCY4HaMX9ocd1MxjYMxa1IeW7HpDcUFj5t3QckLweYFNE
8cQczZ9HrgmNo3EPosF18C67VDF1LBys4nHWSBssD7/VHFCWAOjPKumE7YbpIJee
VjLwlA7CmyzLJiP6q4BRcUZzBX6uQCIKAxM5myMcanDYOqZUhkUIxK5NUR1Dn+Pq
9kAV4inwMidbuJpTUzeplwYBgs8JRZPZZ2fCNKkB4u+Jp9k8aSoa/T6jCRja9OZC
fWeApqzSyG5kFvbrk0ubdTMe1+RSJR8RILbh/UctoX7lv8mbEEEoba9Obi+hODPV
BJct6IWn8sl8F3klAE6uk4azfrWEXgY5LwMBg46Y4mLnJ/YvGWwIOcS+Ko9Apf6y
AiCp4yVZuK5uWi4PbsDoNL9u/u5D2/B5WPXX/ch5z/yJfB004pUexEarC5TKUS7I
yK/jnpwPHBZ1eoLIwRevZFzsO2V3bsElGzWaYK9UaErtiZ4pk5jqJx/fW/LsrOw/
CFVh12UCZ7iahlVGtDl6XeMvH1LqKp22nGs5inVIlzB/FjKMicA049B1g4dcJ/hn
/O+clpahO9OlVN37d+rugthrdecITZMlV3DdYHKY5eUddCBn2NazMIgzqh6rPtN/
qBjvb3npK9vSBWQ+bkxMVHYxSCrfBQuvDFjbZv9WPVmka+sZ42lA+kkmeDWwEtQ7
6Ns31ph2mHugTRMicucsWHgEu1uScAdsfRbAHh/VircrRrcKzOm+wA9ZqC7T9+Il
Kwn7We6oPqzVNZO8Ne3Jg739Iks+UEULvAul6HHEb4wiCr5giTn7qqhPTG1/S0oj
DTUniezD0RJ7KwWosNu/JOxjv+XQevTKZs0A2JkRAmYOOO/EDeVKp2cmX4Kf5nbU
qXtWJYcMsD1EnkQYd9wAtPnSumIDlJ/uG6PEXJYie/USFMcN+pKxKeh/lnkF0mpl
IFFP+ZbyX4qeqqsamP0JrfWdDvPyKX4SLTxECLEtsG51tgRfUAnQ7ZRsNjKD8j+N
uV8x264zI/H2EoXESL1UbjwGE1canWqfNya//Rxkwbf4FQgxrAhMadi6JBUJFrlk
8l31tKLJIxSh/lBSW4nUDrKAfsBJOjeJkOA+ghi3nMT8h2eQXpdjN8Q8/MgwMh9A
Cg6QdRU18k8qXEfn98GQnpE5/A94mQrFxSctrW1VYknnl7L8WB3RmmNYVX2PJzRb
7cTolstwqt7exxUFMmsais793AZPPfGVL++Lk2rNhRiJtmQwlzcR+0UVrsE36U3L
JX6OW8sBuSk+oDTEYbdL7an7SZ8MH+BeHsUxK/ITWeafrOK+Bf5Zm1vzoObjHgKx
yiqy/vIZ1oDd31mz66GYUcQrucHpaPuHFiTU5mUFGL8u5AbRkPp0SdiShmArkuoO
jp129O9vueMAy62nxEYbgK64wc06eThkwx5iG+UGMKBsO6sT1kw9kUNmmeKKkZST
ltNMchjcfdX4ICUt5YcBgiS7M+tv0OF2VGffEdrERJr6ylh+CCgzrkYjoGytUa33
WYv99xB4rs9wE4YazHDdKs3uCspyTIIXJtucsfOol2f24RFgYLETnEsJDQQkMPXw
w0ONUgRY6aGv+XGreg+dWCe+gqCsP8jAIaaAUxyEkuZH7hTHkK5pYfdN/XC8kGdf
Yn4XRlIphy28/HQyIKP/A86igaQ4s2t5J8gK7yh83Lvl3AOE5c/0+u1nSJhuynQB
QmgNaPACOfcFpeQIHACvCELw0L0J3kPqBz917r6nnQz/YL9BLD3HxeSKksxZvs1W
aLc6BpUlbw0nBPz6PKit4Q8y1O/5+lRwAzjrcihqCwDbKCo3hMLYd2Pdj+OZxOcA
0qBhPYdcdybHxsogQN68FzBEThXNIBzn4AUC6ixhTqpeyxElixKq856mttljMLpo
0Vs/02Io/iHogdUvgf3Bt7DBu/X0u8EUklQHCm/UbLc5uCi4Xb0bXkXX6sWL56xB
K9ONjf6x7q2sEYfWZzQYtF9f0ozXAFWFpIydT3P5gQdsxYbY854ZwErf5nKbK157
oX8rLlRJYTrvgMHQd8dkQx2xE4uR19QhNSz6PG+DCcQ2hyxiSfXN/UiZxjuk8NiG
JQ7V6yGG7o1wrs1XSTjK6XExYy97O8Hn8TMr+r2y3bzw3fKgthT6xZuETy1szXXY
R7iO+Lf3NEt+lJVUjwMMzwCuiHow/6x9tkvzwc0TVufyGEsAz9GvujhXmUsemQVN
39B0wZQTN6LIVn0sKts3w5zYlbMdvq7yZKoUNc0sMjCRoqx5T0Jn4LeOy8tSVtZ3
1O7ExAY2FhEMQArzplSOOlRxUURPYTeoDGSUVrxBrlWnkhbeVGuN5yoVYJk+OodC
wBtwZdPT5hfNosQ1AMuyvgFFd9hemYdfKqYMP4QiPBwrcPgK4pbQ71JKnfSnC6nV
jQWKHSj7rHpoV+6/pYkWD7MAuDK58/G3r5VNkFahF5Gub/6NrPU99zwyONkk9W3w
9x2FQY9GkpCUcJHT3DAEa8Oi3y6mndEALxA92z/2Hy9mEwmf1MBo4c45DBHvAL6I
aIZ08gRvSYFL/oMlQlwDnENw3ROTxxBp5LZ8ImNTv0F/xwjNHlHFhcx5XLxEhqwW
UINOvsKlHxRodgn+G6g9bLps6nLOnqDYidn2v/uxwHL9HykRquHHFPkcBgyFeafl
aZs3wRrKyPb+HTE07q3OnkgNkNpL08kAdsRR3PO7vLi+9lI53RCTPqUdipA8iuAI
AztYQ6tOBvxwRez3c8hBlZviQCa40Vt8MtqsLmWpkDxQGy9yh8wNY6IA8CLWAnY4
2F2cFXSVkeSYiR2UdMWN82rKtBbwGO/Jv6AJ5ev5mcU2vfa0/H2KlqFg2/rtwzfL
XcvuyrCJ5O3x6H9Tao3u8gGj/Xo/Jcw+y/rPdWjmD7+wsB/P7Ik07n9b3AzmDdWe
K+J3upgEJ7hO11WHuqor9gRHqlfBbVv1OGK7PwflPa/aXsIZCl1GnkOtecNXgARM
K9u8sjwRXR0H9sPDJp8c2vFROcIP+UVRVgKrLJX4hHgyVH4kXScehSPwbyFwACot
X5ooEm6gpMS90iPRndkzgurJahwtqGult9Hc2/ju45CtVuOOj7uGTYGgoRsek2fK
FK36t5PTSSHREJ9mp9+vTQFZ/b0cEzIr+pvf2nG88MeiMf2JF4CMTS1sDQO1Hbqf
6vrqw1CYxTuZIfcFbMRJgnWlrhBOkirxAoeAOwDcEc89v2cEtIvFDh3IlbjpZ//+
13R/k/I4f6FSl5wQZV53Peezm0au3jBgRiFKd0J1lIVe4AJ4St+4coerlT0gXwFu
tcQykcK4P2O7UCWGHa31oNZspCGbeoktwuxfhmp34NAj3fwsEupXrTxqNUTdAdOc
TqlknD8ka7mWqj4gF0KEs7YxlUTiE6rCvSYnZ0x3ok77ki/IDCH0FPISDc0GlcrU
+bPxCUYWaHmpu9Q1t7UY+uTj7CanMvBDxF9sGW8sfRtZUbYXBQ3VI/PyTrAtekwy
o2nfQViVyH6TFezos87V4+De9f6KaZEsRk7HOsbMbYbbWqTKXerhXZwXN+dokx8m
EGElP3D9KxiQAiNVkWdVTS8yi2EuxL9iGAkJd/GNkQVFLfaisRYcGYxIeOdln7DH
fOiUXN/4J68JVaKJmy5Td5MipySFu89THXJyC53z66wzPkFdk/cxf8zMfpo0JcyD
9xTh7M6Knrd3LrM3TU2J1MzymaeRbDDzKp6t3T4OKu8h766Gfn6lNTAST8XQ7wJy
6mXnFP8IdwjHGGDLz8GPNll5ro1g7ByPd2oYkFiDJ2QfjTdibeZ6bXbHwaZ14pfz
hRYqFbwEJmLoaaUAGsVAQzjxTQTmv1hFRecsjZLaG6T0CQIVGn6HeAwBuxISTP8A
/WHy6MD0481wp6gDf/L8DN5gYOVhQIcWuE37oTgBiciUnGXOBT+ZM6tIUtO35RWE
mCMIFis4hDAJGmP1qmLL6h3PVFHAof8myWhOD7gjRuiRBNyrTApiXoGITo+m/HCE
+5KeL2Mv+n3/R4tZ2htsNrHyDp+9TbHSZy9OOerpVLpYdDoM7HvrmyAzKQp+g/p5
vckd5xopCZSX8bx3BFCEt2jabnaPPmj8XGSsGZLeePhfpglNQRYgn6qulv3OrhLE
pCGANzIdwxh4nL2wKBgcMpKImjEM02eg3OGhzxnKKEZ5VOZpLYNuSEpcR9Q/Z8AW
XE9IhWw1L+blnDWZdM3LylnQpzcFt5w0DAJhpTfZJmKgMMIfOtlZAfQhR294Gq9E
DxI89pTHX2Hq0Ami5UzNTZ20bgTIrzjZjxFWemHpB0zmrJMgwYrbJRtkrmBRQJNX
4TRESrNdP5Ery14sRE2RmWPbh25C3ZDFykiw9lHzVyKyVgJ4l8Jb+6FA7BT6pM04
ljwmOEnx0fuFTkHz3NLPiLACEV3R3v9nhPFQLE/Lwc7oKQ1iBjWt3+N7HZBQdylC
S/TCNPrDy1GZ1R/mc1W67Z+EYEybEAAYob7q1f/UuNfqLIepZHWhzKIpKpME62nz
WPqvARo16IkYd/tJoKnncBlSTpAjrZe/TRnt7+IqkZC0qdIvAAMEg9afOO5gwD7Q
fJshcIPqoxLFksUa+w2n7ifHnNOeU1qfxugp5DLCpZyQDQe7j1I97Mc86SsGn7SF
3nd2v+uwseIyzUfy9EO//0WZuGyvcAFxx1hQqgJo+9e7pmC3RxDwTgoee09nUYLS
wVFfFVUzH0xsKG7uOcP6yKGCcb9rUYnWqJzfFTMgM1k1V5ahSAQPSCyhkh6pYRkA
0oyRfgjojnwZ4Kb6B+b02/I84Dplw6PtVO9fcPvKEghtWZ8RBfMPjBSFe/V1KBKi
NPtdafg8JP0Dbks4xuDtmjCzI1T8mGZgavJbxSRPc1dTxoCP8d7+lgD+WpbMLqY2
xyIFYBt5kEVMTUN4chYTq1pPHWjK/6EFTFPoCORt2fd7vnNkk7iYYi29Trl8v6RK
8S8wlTAn+OTJNedmXV1B2gLzO476Y411aFua+prYbnJfFwG06rmk7HmdV8t8mHE5
vFDKwoVosD9/LQc03geIfyuDV8ubA4TXHly/RpEsCkA17INpVC9zau0ZP6nbIEFF
PdU2W4w6wg45EK8BCjk4pLPScvqczeXeapPg0HQgWbKqNXQ3v97lGTjn0BM+qpct

//pragma protect end_data_block
//pragma protect digest_block
MeaHDqM2BRv+XIQTTNbelE46pDU=
//pragma protect end_digest_block
//pragma protect end_protected
